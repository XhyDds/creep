module priv (
    output [1:0]PLV
);
    
endmodule