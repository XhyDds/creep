module data_pre#(

)(

);
endmodule