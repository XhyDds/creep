module SUC ( //强序非缓存刷新pc
    input      clk,
    input      rstn,
    
);
    
endmodule //SUC
