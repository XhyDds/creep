module priv (
    
);
    
endmodule