module ReturnBuffer #(
    parameter   index_width=4,
                offset_width=2,
) (
    input   wire    clk,
    input   wire    rst,
    
);
    
endmodule