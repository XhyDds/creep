module priv (
    output [1:0]PLV
);
    assign PLV=0;
endmodule
