
`timescale 1ns / 1ps
module cache_tb();

localparam INDEX_WIDTH          = 2;
localparam WORD_OFFSET_WIDTH    = 2;
localparam TOTAL_WORD_NUM       = 1024;

// cache test
reg [31:0]  i_addr_rom [TOTAL_WORD_NUM];
reg [31:0]  d_addr_rom [TOTAL_WORD_NUM];
reg [31:0]  data_ram [TOTAL_WORD_NUM];
reg         wvalid_rom [TOTAL_WORD_NUM];
reg [31:0]  wdata_rom [TOTAL_WORD_NUM];
reg [31:0]  i_test_index = 0;
reg [31:0]  d_test_index = 0;
reg clk = 1'b1, rstn = 1'b0;

initial #5 rstn = 1'b1; 
always #1 clk = ~clk;

// generate data_ram
initial begin
    data_ram[    0] = 'h00000000; 	    data_ram[    1] = 'h00000001; 	    data_ram[    2] = 'h00000002; 	    data_ram[    3] = 'h00000003; 	    data_ram[    4] = 'h00000004; 	    data_ram[    5] = 'h00000005; 	    data_ram[    6] = 'h00000006; 	    data_ram[    7] = 'h00000007; 	
    data_ram[    8] = 'h00000008; 	    data_ram[    9] = 'h00000009; 	    data_ram[   10] = 'h0000000a; 	    data_ram[   11] = 'h0000000b; 	    data_ram[   12] = 'h0000000c; 	    data_ram[   13] = 'h0000000d; 	    data_ram[   14] = 'h0000000e; 	    data_ram[   15] = 'h0000000f; 	
    data_ram[   16] = 'h00000010; 	    data_ram[   17] = 'h00000011; 	    data_ram[   18] = 'h00000012; 	    data_ram[   19] = 'h00000013; 	    data_ram[   20] = 'h00000014; 	    data_ram[   21] = 'h00000015; 	    data_ram[   22] = 'h00000016; 	    data_ram[   23] = 'h00000017; 	
    data_ram[   24] = 'h00000018; 	    data_ram[   25] = 'h00000019; 	    data_ram[   26] = 'h0000001a; 	    data_ram[   27] = 'h0000001b; 	    data_ram[   28] = 'h0000001c; 	    data_ram[   29] = 'h0000001d; 	    data_ram[   30] = 'h0000001e; 	    data_ram[   31] = 'h0000001f; 	
    data_ram[   32] = 'h00000020; 	    data_ram[   33] = 'h00000021; 	    data_ram[   34] = 'h00000022; 	    data_ram[   35] = 'h00000023; 	    data_ram[   36] = 'h00000024; 	    data_ram[   37] = 'h00000025; 	    data_ram[   38] = 'h00000026; 	    data_ram[   39] = 'h00000027; 	
    data_ram[   40] = 'h00000028; 	    data_ram[   41] = 'h00000029; 	    data_ram[   42] = 'h0000002a; 	    data_ram[   43] = 'h0000002b; 	    data_ram[   44] = 'h0000002c; 	    data_ram[   45] = 'h0000002d; 	    data_ram[   46] = 'h0000002e; 	    data_ram[   47] = 'h0000002f; 	
    data_ram[   48] = 'h00000030; 	    data_ram[   49] = 'h00000031; 	    data_ram[   50] = 'h00000032; 	    data_ram[   51] = 'h00000033; 	    data_ram[   52] = 'h00000034; 	    data_ram[   53] = 'h00000035; 	    data_ram[   54] = 'h00000036; 	    data_ram[   55] = 'h00000037; 	
    data_ram[   56] = 'h00000038; 	    data_ram[   57] = 'h00000039; 	    data_ram[   58] = 'h0000003a; 	    data_ram[   59] = 'h0000003b; 	    data_ram[   60] = 'h0000003c; 	    data_ram[   61] = 'h0000003d; 	    data_ram[   62] = 'h0000003e; 	    data_ram[   63] = 'h0000003f; 	
    data_ram[   64] = 'h00000040; 	    data_ram[   65] = 'h00000041; 	    data_ram[   66] = 'h00000042; 	    data_ram[   67] = 'h00000043; 	    data_ram[   68] = 'h00000044; 	    data_ram[   69] = 'h00000045; 	    data_ram[   70] = 'h00000046; 	    data_ram[   71] = 'h00000047; 	
    data_ram[   72] = 'h00000048; 	    data_ram[   73] = 'h00000049; 	    data_ram[   74] = 'h0000004a; 	    data_ram[   75] = 'h0000004b; 	    data_ram[   76] = 'h0000004c; 	    data_ram[   77] = 'h0000004d; 	    data_ram[   78] = 'h0000004e; 	    data_ram[   79] = 'h0000004f; 	
    data_ram[   80] = 'h00000050; 	    data_ram[   81] = 'h00000051; 	    data_ram[   82] = 'h00000052; 	    data_ram[   83] = 'h00000053; 	    data_ram[   84] = 'h00000054; 	    data_ram[   85] = 'h00000055; 	    data_ram[   86] = 'h00000056; 	    data_ram[   87] = 'h00000057; 	
    data_ram[   88] = 'h00000058; 	    data_ram[   89] = 'h00000059; 	    data_ram[   90] = 'h0000005a; 	    data_ram[   91] = 'h0000005b; 	    data_ram[   92] = 'h0000005c; 	    data_ram[   93] = 'h0000005d; 	    data_ram[   94] = 'h0000005e; 	    data_ram[   95] = 'h0000005f; 	
    data_ram[   96] = 'h00000060; 	    data_ram[   97] = 'h00000061; 	    data_ram[   98] = 'h00000062; 	    data_ram[   99] = 'h00000063; 	    data_ram[  100] = 'h00000064; 	    data_ram[  101] = 'h00000065; 	    data_ram[  102] = 'h00000066; 	    data_ram[  103] = 'h00000067; 	
    data_ram[  104] = 'h00000068; 	    data_ram[  105] = 'h00000069; 	    data_ram[  106] = 'h0000006a; 	    data_ram[  107] = 'h0000006b; 	    data_ram[  108] = 'h0000006c; 	    data_ram[  109] = 'h0000006d; 	    data_ram[  110] = 'h0000006e; 	    data_ram[  111] = 'h0000006f; 	
    data_ram[  112] = 'h00000070; 	    data_ram[  113] = 'h00000071; 	    data_ram[  114] = 'h00000072; 	    data_ram[  115] = 'h00000073; 	    data_ram[  116] = 'h00000074; 	    data_ram[  117] = 'h00000075; 	    data_ram[  118] = 'h00000076; 	    data_ram[  119] = 'h00000077; 	
    data_ram[  120] = 'h00000078; 	    data_ram[  121] = 'h00000079; 	    data_ram[  122] = 'h0000007a; 	    data_ram[  123] = 'h0000007b; 	    data_ram[  124] = 'h0000007c; 	    data_ram[  125] = 'h0000007d; 	    data_ram[  126] = 'h0000007e; 	    data_ram[  127] = 'h0000007f; 	
    data_ram[  128] = 'h00000080; 	    data_ram[  129] = 'h00000081; 	    data_ram[  130] = 'h00000082; 	    data_ram[  131] = 'h00000083; 	    data_ram[  132] = 'h00000084; 	    data_ram[  133] = 'h00000085; 	    data_ram[  134] = 'h00000086; 	    data_ram[  135] = 'h00000087; 	
    data_ram[  136] = 'h00000088; 	    data_ram[  137] = 'h00000089; 	    data_ram[  138] = 'h0000008a; 	    data_ram[  139] = 'h0000008b; 	    data_ram[  140] = 'h0000008c; 	    data_ram[  141] = 'h0000008d; 	    data_ram[  142] = 'h0000008e; 	    data_ram[  143] = 'h0000008f; 	
    data_ram[  144] = 'h00000090; 	    data_ram[  145] = 'h00000091; 	    data_ram[  146] = 'h00000092; 	    data_ram[  147] = 'h00000093; 	    data_ram[  148] = 'h00000094; 	    data_ram[  149] = 'h00000095; 	    data_ram[  150] = 'h00000096; 	    data_ram[  151] = 'h00000097; 	
    data_ram[  152] = 'h00000098; 	    data_ram[  153] = 'h00000099; 	    data_ram[  154] = 'h0000009a; 	    data_ram[  155] = 'h0000009b; 	    data_ram[  156] = 'h0000009c; 	    data_ram[  157] = 'h0000009d; 	    data_ram[  158] = 'h0000009e; 	    data_ram[  159] = 'h0000009f; 	
    data_ram[  160] = 'h000000a0; 	    data_ram[  161] = 'h000000a1; 	    data_ram[  162] = 'h000000a2; 	    data_ram[  163] = 'h000000a3; 	    data_ram[  164] = 'h000000a4; 	    data_ram[  165] = 'h000000a5; 	    data_ram[  166] = 'h000000a6; 	    data_ram[  167] = 'h000000a7; 	
    data_ram[  168] = 'h000000a8; 	    data_ram[  169] = 'h000000a9; 	    data_ram[  170] = 'h000000aa; 	    data_ram[  171] = 'h000000ab; 	    data_ram[  172] = 'h000000ac; 	    data_ram[  173] = 'h000000ad; 	    data_ram[  174] = 'h000000ae; 	    data_ram[  175] = 'h000000af; 	
    data_ram[  176] = 'h000000b0; 	    data_ram[  177] = 'h000000b1; 	    data_ram[  178] = 'h000000b2; 	    data_ram[  179] = 'h000000b3; 	    data_ram[  180] = 'h000000b4; 	    data_ram[  181] = 'h000000b5; 	    data_ram[  182] = 'h000000b6; 	    data_ram[  183] = 'h000000b7; 	
    data_ram[  184] = 'h000000b8; 	    data_ram[  185] = 'h000000b9; 	    data_ram[  186] = 'h000000ba; 	    data_ram[  187] = 'h000000bb; 	    data_ram[  188] = 'h000000bc; 	    data_ram[  189] = 'h000000bd; 	    data_ram[  190] = 'h000000be; 	    data_ram[  191] = 'h000000bf; 	
    data_ram[  192] = 'h000000c0; 	    data_ram[  193] = 'h000000c1; 	    data_ram[  194] = 'h000000c2; 	    data_ram[  195] = 'h000000c3; 	    data_ram[  196] = 'h000000c4; 	    data_ram[  197] = 'h000000c5; 	    data_ram[  198] = 'h000000c6; 	    data_ram[  199] = 'h000000c7; 	
    data_ram[  200] = 'h000000c8; 	    data_ram[  201] = 'h000000c9; 	    data_ram[  202] = 'h000000ca; 	    data_ram[  203] = 'h000000cb; 	    data_ram[  204] = 'h000000cc; 	    data_ram[  205] = 'h000000cd; 	    data_ram[  206] = 'h000000ce; 	    data_ram[  207] = 'h000000cf; 	
    data_ram[  208] = 'h000000d0; 	    data_ram[  209] = 'h000000d1; 	    data_ram[  210] = 'h000000d2; 	    data_ram[  211] = 'h000000d3; 	    data_ram[  212] = 'h000000d4; 	    data_ram[  213] = 'h000000d5; 	    data_ram[  214] = 'h000000d6; 	    data_ram[  215] = 'h000000d7; 	
    data_ram[  216] = 'h000000d8; 	    data_ram[  217] = 'h000000d9; 	    data_ram[  218] = 'h000000da; 	    data_ram[  219] = 'h000000db; 	    data_ram[  220] = 'h000000dc; 	    data_ram[  221] = 'h000000dd; 	    data_ram[  222] = 'h000000de; 	    data_ram[  223] = 'h000000df; 	
    data_ram[  224] = 'h000000e0; 	    data_ram[  225] = 'h000000e1; 	    data_ram[  226] = 'h000000e2; 	    data_ram[  227] = 'h000000e3; 	    data_ram[  228] = 'h000000e4; 	    data_ram[  229] = 'h000000e5; 	    data_ram[  230] = 'h000000e6; 	    data_ram[  231] = 'h000000e7; 	
    data_ram[  232] = 'h000000e8; 	    data_ram[  233] = 'h000000e9; 	    data_ram[  234] = 'h000000ea; 	    data_ram[  235] = 'h000000eb; 	    data_ram[  236] = 'h000000ec; 	    data_ram[  237] = 'h000000ed; 	    data_ram[  238] = 'h000000ee; 	    data_ram[  239] = 'h000000ef; 	
    data_ram[  240] = 'h000000f0; 	    data_ram[  241] = 'h000000f1; 	    data_ram[  242] = 'h000000f2; 	    data_ram[  243] = 'h000000f3; 	    data_ram[  244] = 'h000000f4; 	    data_ram[  245] = 'h000000f5; 	    data_ram[  246] = 'h000000f6; 	    data_ram[  247] = 'h000000f7; 	
    data_ram[  248] = 'h000000f8; 	    data_ram[  249] = 'h000000f9; 	    data_ram[  250] = 'h000000fa; 	    data_ram[  251] = 'h000000fb; 	    data_ram[  252] = 'h000000fc; 	    data_ram[  253] = 'h000000fd; 	    data_ram[  254] = 'h000000fe; 	    data_ram[  255] = 'h000000ff; 	
    data_ram[  256] = 'h00000100; 	    data_ram[  257] = 'h00000101; 	    data_ram[  258] = 'h00000102; 	    data_ram[  259] = 'h00000103; 	    data_ram[  260] = 'h00000104; 	    data_ram[  261] = 'h00000105; 	    data_ram[  262] = 'h00000106; 	    data_ram[  263] = 'h00000107; 	
    data_ram[  264] = 'h00000108; 	    data_ram[  265] = 'h00000109; 	    data_ram[  266] = 'h0000010a; 	    data_ram[  267] = 'h0000010b; 	    data_ram[  268] = 'h0000010c; 	    data_ram[  269] = 'h0000010d; 	    data_ram[  270] = 'h0000010e; 	    data_ram[  271] = 'h0000010f; 	
    data_ram[  272] = 'h00000110; 	    data_ram[  273] = 'h00000111; 	    data_ram[  274] = 'h00000112; 	    data_ram[  275] = 'h00000113; 	    data_ram[  276] = 'h00000114; 	    data_ram[  277] = 'h00000115; 	    data_ram[  278] = 'h00000116; 	    data_ram[  279] = 'h00000117; 	
    data_ram[  280] = 'h00000118; 	    data_ram[  281] = 'h00000119; 	    data_ram[  282] = 'h0000011a; 	    data_ram[  283] = 'h0000011b; 	    data_ram[  284] = 'h0000011c; 	    data_ram[  285] = 'h0000011d; 	    data_ram[  286] = 'h0000011e; 	    data_ram[  287] = 'h0000011f; 	
    data_ram[  288] = 'h00000120; 	    data_ram[  289] = 'h00000121; 	    data_ram[  290] = 'h00000122; 	    data_ram[  291] = 'h00000123; 	    data_ram[  292] = 'h00000124; 	    data_ram[  293] = 'h00000125; 	    data_ram[  294] = 'h00000126; 	    data_ram[  295] = 'h00000127; 	
    data_ram[  296] = 'h00000128; 	    data_ram[  297] = 'h00000129; 	    data_ram[  298] = 'h0000012a; 	    data_ram[  299] = 'h0000012b; 	    data_ram[  300] = 'h0000012c; 	    data_ram[  301] = 'h0000012d; 	    data_ram[  302] = 'h0000012e; 	    data_ram[  303] = 'h0000012f; 	
    data_ram[  304] = 'h00000130; 	    data_ram[  305] = 'h00000131; 	    data_ram[  306] = 'h00000132; 	    data_ram[  307] = 'h00000133; 	    data_ram[  308] = 'h00000134; 	    data_ram[  309] = 'h00000135; 	    data_ram[  310] = 'h00000136; 	    data_ram[  311] = 'h00000137; 	
    data_ram[  312] = 'h00000138; 	    data_ram[  313] = 'h00000139; 	    data_ram[  314] = 'h0000013a; 	    data_ram[  315] = 'h0000013b; 	    data_ram[  316] = 'h0000013c; 	    data_ram[  317] = 'h0000013d; 	    data_ram[  318] = 'h0000013e; 	    data_ram[  319] = 'h0000013f; 	
    data_ram[  320] = 'h00000140; 	    data_ram[  321] = 'h00000141; 	    data_ram[  322] = 'h00000142; 	    data_ram[  323] = 'h00000143; 	    data_ram[  324] = 'h00000144; 	    data_ram[  325] = 'h00000145; 	    data_ram[  326] = 'h00000146; 	    data_ram[  327] = 'h00000147; 	
    data_ram[  328] = 'h00000148; 	    data_ram[  329] = 'h00000149; 	    data_ram[  330] = 'h0000014a; 	    data_ram[  331] = 'h0000014b; 	    data_ram[  332] = 'h0000014c; 	    data_ram[  333] = 'h0000014d; 	    data_ram[  334] = 'h0000014e; 	    data_ram[  335] = 'h0000014f; 	
    data_ram[  336] = 'h00000150; 	    data_ram[  337] = 'h00000151; 	    data_ram[  338] = 'h00000152; 	    data_ram[  339] = 'h00000153; 	    data_ram[  340] = 'h00000154; 	    data_ram[  341] = 'h00000155; 	    data_ram[  342] = 'h00000156; 	    data_ram[  343] = 'h00000157; 	
    data_ram[  344] = 'h00000158; 	    data_ram[  345] = 'h00000159; 	    data_ram[  346] = 'h0000015a; 	    data_ram[  347] = 'h0000015b; 	    data_ram[  348] = 'h0000015c; 	    data_ram[  349] = 'h0000015d; 	    data_ram[  350] = 'h0000015e; 	    data_ram[  351] = 'h0000015f; 	
    data_ram[  352] = 'h00000160; 	    data_ram[  353] = 'h00000161; 	    data_ram[  354] = 'h00000162; 	    data_ram[  355] = 'h00000163; 	    data_ram[  356] = 'h00000164; 	    data_ram[  357] = 'h00000165; 	    data_ram[  358] = 'h00000166; 	    data_ram[  359] = 'h00000167; 	
    data_ram[  360] = 'h00000168; 	    data_ram[  361] = 'h00000169; 	    data_ram[  362] = 'h0000016a; 	    data_ram[  363] = 'h0000016b; 	    data_ram[  364] = 'h0000016c; 	    data_ram[  365] = 'h0000016d; 	    data_ram[  366] = 'h0000016e; 	    data_ram[  367] = 'h0000016f; 	
    data_ram[  368] = 'h00000170; 	    data_ram[  369] = 'h00000171; 	    data_ram[  370] = 'h00000172; 	    data_ram[  371] = 'h00000173; 	    data_ram[  372] = 'h00000174; 	    data_ram[  373] = 'h00000175; 	    data_ram[  374] = 'h00000176; 	    data_ram[  375] = 'h00000177; 	
    data_ram[  376] = 'h00000178; 	    data_ram[  377] = 'h00000179; 	    data_ram[  378] = 'h0000017a; 	    data_ram[  379] = 'h0000017b; 	    data_ram[  380] = 'h0000017c; 	    data_ram[  381] = 'h0000017d; 	    data_ram[  382] = 'h0000017e; 	    data_ram[  383] = 'h0000017f; 	
    data_ram[  384] = 'h00000180; 	    data_ram[  385] = 'h00000181; 	    data_ram[  386] = 'h00000182; 	    data_ram[  387] = 'h00000183; 	    data_ram[  388] = 'h00000184; 	    data_ram[  389] = 'h00000185; 	    data_ram[  390] = 'h00000186; 	    data_ram[  391] = 'h00000187; 	
    data_ram[  392] = 'h00000188; 	    data_ram[  393] = 'h00000189; 	    data_ram[  394] = 'h0000018a; 	    data_ram[  395] = 'h0000018b; 	    data_ram[  396] = 'h0000018c; 	    data_ram[  397] = 'h0000018d; 	    data_ram[  398] = 'h0000018e; 	    data_ram[  399] = 'h0000018f; 	
    data_ram[  400] = 'h00000190; 	    data_ram[  401] = 'h00000191; 	    data_ram[  402] = 'h00000192; 	    data_ram[  403] = 'h00000193; 	    data_ram[  404] = 'h00000194; 	    data_ram[  405] = 'h00000195; 	    data_ram[  406] = 'h00000196; 	    data_ram[  407] = 'h00000197; 	
    data_ram[  408] = 'h00000198; 	    data_ram[  409] = 'h00000199; 	    data_ram[  410] = 'h0000019a; 	    data_ram[  411] = 'h0000019b; 	    data_ram[  412] = 'h0000019c; 	    data_ram[  413] = 'h0000019d; 	    data_ram[  414] = 'h0000019e; 	    data_ram[  415] = 'h0000019f; 	
    data_ram[  416] = 'h000001a0; 	    data_ram[  417] = 'h000001a1; 	    data_ram[  418] = 'h000001a2; 	    data_ram[  419] = 'h000001a3; 	    data_ram[  420] = 'h000001a4; 	    data_ram[  421] = 'h000001a5; 	    data_ram[  422] = 'h000001a6; 	    data_ram[  423] = 'h000001a7; 	
    data_ram[  424] = 'h000001a8; 	    data_ram[  425] = 'h000001a9; 	    data_ram[  426] = 'h000001aa; 	    data_ram[  427] = 'h000001ab; 	    data_ram[  428] = 'h000001ac; 	    data_ram[  429] = 'h000001ad; 	    data_ram[  430] = 'h000001ae; 	    data_ram[  431] = 'h000001af; 	
    data_ram[  432] = 'h000001b0; 	    data_ram[  433] = 'h000001b1; 	    data_ram[  434] = 'h000001b2; 	    data_ram[  435] = 'h000001b3; 	    data_ram[  436] = 'h000001b4; 	    data_ram[  437] = 'h000001b5; 	    data_ram[  438] = 'h000001b6; 	    data_ram[  439] = 'h000001b7; 	
    data_ram[  440] = 'h000001b8; 	    data_ram[  441] = 'h000001b9; 	    data_ram[  442] = 'h000001ba; 	    data_ram[  443] = 'h000001bb; 	    data_ram[  444] = 'h000001bc; 	    data_ram[  445] = 'h000001bd; 	    data_ram[  446] = 'h000001be; 	    data_ram[  447] = 'h000001bf; 	
    data_ram[  448] = 'h000001c0; 	    data_ram[  449] = 'h000001c1; 	    data_ram[  450] = 'h000001c2; 	    data_ram[  451] = 'h000001c3; 	    data_ram[  452] = 'h000001c4; 	    data_ram[  453] = 'h000001c5; 	    data_ram[  454] = 'h000001c6; 	    data_ram[  455] = 'h000001c7; 	
    data_ram[  456] = 'h000001c8; 	    data_ram[  457] = 'h000001c9; 	    data_ram[  458] = 'h000001ca; 	    data_ram[  459] = 'h000001cb; 	    data_ram[  460] = 'h000001cc; 	    data_ram[  461] = 'h000001cd; 	    data_ram[  462] = 'h000001ce; 	    data_ram[  463] = 'h000001cf; 	
    data_ram[  464] = 'h000001d0; 	    data_ram[  465] = 'h000001d1; 	    data_ram[  466] = 'h000001d2; 	    data_ram[  467] = 'h000001d3; 	    data_ram[  468] = 'h000001d4; 	    data_ram[  469] = 'h000001d5; 	    data_ram[  470] = 'h000001d6; 	    data_ram[  471] = 'h000001d7; 	
    data_ram[  472] = 'h000001d8; 	    data_ram[  473] = 'h000001d9; 	    data_ram[  474] = 'h000001da; 	    data_ram[  475] = 'h000001db; 	    data_ram[  476] = 'h000001dc; 	    data_ram[  477] = 'h000001dd; 	    data_ram[  478] = 'h000001de; 	    data_ram[  479] = 'h000001df; 	
    data_ram[  480] = 'h000001e0; 	    data_ram[  481] = 'h000001e1; 	    data_ram[  482] = 'h000001e2; 	    data_ram[  483] = 'h000001e3; 	    data_ram[  484] = 'h000001e4; 	    data_ram[  485] = 'h000001e5; 	    data_ram[  486] = 'h000001e6; 	    data_ram[  487] = 'h000001e7; 	
    data_ram[  488] = 'h000001e8; 	    data_ram[  489] = 'h000001e9; 	    data_ram[  490] = 'h000001ea; 	    data_ram[  491] = 'h000001eb; 	    data_ram[  492] = 'h000001ec; 	    data_ram[  493] = 'h000001ed; 	    data_ram[  494] = 'h000001ee; 	    data_ram[  495] = 'h000001ef; 	
    data_ram[  496] = 'h000001f0; 	    data_ram[  497] = 'h000001f1; 	    data_ram[  498] = 'h000001f2; 	    data_ram[  499] = 'h000001f3; 	    data_ram[  500] = 'h000001f4; 	    data_ram[  501] = 'h000001f5; 	    data_ram[  502] = 'h000001f6; 	    data_ram[  503] = 'h000001f7; 	
    data_ram[  504] = 'h000001f8; 	    data_ram[  505] = 'h000001f9; 	    data_ram[  506] = 'h000001fa; 	    data_ram[  507] = 'h000001fb; 	    data_ram[  508] = 'h000001fc; 	    data_ram[  509] = 'h000001fd; 	    data_ram[  510] = 'h000001fe; 	    data_ram[  511] = 'h000001ff; 	
    data_ram[  512] = 'h00000200; 	    data_ram[  513] = 'h00000201; 	    data_ram[  514] = 'h00000202; 	    data_ram[  515] = 'h00000203; 	    data_ram[  516] = 'h00000204; 	    data_ram[  517] = 'h00000205; 	    data_ram[  518] = 'h00000206; 	    data_ram[  519] = 'h00000207; 	
    data_ram[  520] = 'h00000208; 	    data_ram[  521] = 'h00000209; 	    data_ram[  522] = 'h0000020a; 	    data_ram[  523] = 'h0000020b; 	    data_ram[  524] = 'h0000020c; 	    data_ram[  525] = 'h0000020d; 	    data_ram[  526] = 'h0000020e; 	    data_ram[  527] = 'h0000020f; 	
    data_ram[  528] = 'h00000210; 	    data_ram[  529] = 'h00000211; 	    data_ram[  530] = 'h00000212; 	    data_ram[  531] = 'h00000213; 	    data_ram[  532] = 'h00000214; 	    data_ram[  533] = 'h00000215; 	    data_ram[  534] = 'h00000216; 	    data_ram[  535] = 'h00000217; 	
    data_ram[  536] = 'h00000218; 	    data_ram[  537] = 'h00000219; 	    data_ram[  538] = 'h0000021a; 	    data_ram[  539] = 'h0000021b; 	    data_ram[  540] = 'h0000021c; 	    data_ram[  541] = 'h0000021d; 	    data_ram[  542] = 'h0000021e; 	    data_ram[  543] = 'h0000021f; 	
    data_ram[  544] = 'h00000220; 	    data_ram[  545] = 'h00000221; 	    data_ram[  546] = 'h00000222; 	    data_ram[  547] = 'h00000223; 	    data_ram[  548] = 'h00000224; 	    data_ram[  549] = 'h00000225; 	    data_ram[  550] = 'h00000226; 	    data_ram[  551] = 'h00000227; 	
    data_ram[  552] = 'h00000228; 	    data_ram[  553] = 'h00000229; 	    data_ram[  554] = 'h0000022a; 	    data_ram[  555] = 'h0000022b; 	    data_ram[  556] = 'h0000022c; 	    data_ram[  557] = 'h0000022d; 	    data_ram[  558] = 'h0000022e; 	    data_ram[  559] = 'h0000022f; 	
    data_ram[  560] = 'h00000230; 	    data_ram[  561] = 'h00000231; 	    data_ram[  562] = 'h00000232; 	    data_ram[  563] = 'h00000233; 	    data_ram[  564] = 'h00000234; 	    data_ram[  565] = 'h00000235; 	    data_ram[  566] = 'h00000236; 	    data_ram[  567] = 'h00000237; 	
    data_ram[  568] = 'h00000238; 	    data_ram[  569] = 'h00000239; 	    data_ram[  570] = 'h0000023a; 	    data_ram[  571] = 'h0000023b; 	    data_ram[  572] = 'h0000023c; 	    data_ram[  573] = 'h0000023d; 	    data_ram[  574] = 'h0000023e; 	    data_ram[  575] = 'h0000023f; 	
    data_ram[  576] = 'h00000240; 	    data_ram[  577] = 'h00000241; 	    data_ram[  578] = 'h00000242; 	    data_ram[  579] = 'h00000243; 	    data_ram[  580] = 'h00000244; 	    data_ram[  581] = 'h00000245; 	    data_ram[  582] = 'h00000246; 	    data_ram[  583] = 'h00000247; 	
    data_ram[  584] = 'h00000248; 	    data_ram[  585] = 'h00000249; 	    data_ram[  586] = 'h0000024a; 	    data_ram[  587] = 'h0000024b; 	    data_ram[  588] = 'h0000024c; 	    data_ram[  589] = 'h0000024d; 	    data_ram[  590] = 'h0000024e; 	    data_ram[  591] = 'h0000024f; 	
    data_ram[  592] = 'h00000250; 	    data_ram[  593] = 'h00000251; 	    data_ram[  594] = 'h00000252; 	    data_ram[  595] = 'h00000253; 	    data_ram[  596] = 'h00000254; 	    data_ram[  597] = 'h00000255; 	    data_ram[  598] = 'h00000256; 	    data_ram[  599] = 'h00000257; 	
    data_ram[  600] = 'h00000258; 	    data_ram[  601] = 'h00000259; 	    data_ram[  602] = 'h0000025a; 	    data_ram[  603] = 'h0000025b; 	    data_ram[  604] = 'h0000025c; 	    data_ram[  605] = 'h0000025d; 	    data_ram[  606] = 'h0000025e; 	    data_ram[  607] = 'h0000025f; 	
    data_ram[  608] = 'h00000260; 	    data_ram[  609] = 'h00000261; 	    data_ram[  610] = 'h00000262; 	    data_ram[  611] = 'h00000263; 	    data_ram[  612] = 'h00000264; 	    data_ram[  613] = 'h00000265; 	    data_ram[  614] = 'h00000266; 	    data_ram[  615] = 'h00000267; 	
    data_ram[  616] = 'h00000268; 	    data_ram[  617] = 'h00000269; 	    data_ram[  618] = 'h0000026a; 	    data_ram[  619] = 'h0000026b; 	    data_ram[  620] = 'h0000026c; 	    data_ram[  621] = 'h0000026d; 	    data_ram[  622] = 'h0000026e; 	    data_ram[  623] = 'h0000026f; 	
    data_ram[  624] = 'h00000270; 	    data_ram[  625] = 'h00000271; 	    data_ram[  626] = 'h00000272; 	    data_ram[  627] = 'h00000273; 	    data_ram[  628] = 'h00000274; 	    data_ram[  629] = 'h00000275; 	    data_ram[  630] = 'h00000276; 	    data_ram[  631] = 'h00000277; 	
    data_ram[  632] = 'h00000278; 	    data_ram[  633] = 'h00000279; 	    data_ram[  634] = 'h0000027a; 	    data_ram[  635] = 'h0000027b; 	    data_ram[  636] = 'h0000027c; 	    data_ram[  637] = 'h0000027d; 	    data_ram[  638] = 'h0000027e; 	    data_ram[  639] = 'h0000027f; 	
    data_ram[  640] = 'h00000280; 	    data_ram[  641] = 'h00000281; 	    data_ram[  642] = 'h00000282; 	    data_ram[  643] = 'h00000283; 	    data_ram[  644] = 'h00000284; 	    data_ram[  645] = 'h00000285; 	    data_ram[  646] = 'h00000286; 	    data_ram[  647] = 'h00000287; 	
    data_ram[  648] = 'h00000288; 	    data_ram[  649] = 'h00000289; 	    data_ram[  650] = 'h0000028a; 	    data_ram[  651] = 'h0000028b; 	    data_ram[  652] = 'h0000028c; 	    data_ram[  653] = 'h0000028d; 	    data_ram[  654] = 'h0000028e; 	    data_ram[  655] = 'h0000028f; 	
    data_ram[  656] = 'h00000290; 	    data_ram[  657] = 'h00000291; 	    data_ram[  658] = 'h00000292; 	    data_ram[  659] = 'h00000293; 	    data_ram[  660] = 'h00000294; 	    data_ram[  661] = 'h00000295; 	    data_ram[  662] = 'h00000296; 	    data_ram[  663] = 'h00000297; 	
    data_ram[  664] = 'h00000298; 	    data_ram[  665] = 'h00000299; 	    data_ram[  666] = 'h0000029a; 	    data_ram[  667] = 'h0000029b; 	    data_ram[  668] = 'h0000029c; 	    data_ram[  669] = 'h0000029d; 	    data_ram[  670] = 'h0000029e; 	    data_ram[  671] = 'h0000029f; 	
    data_ram[  672] = 'h000002a0; 	    data_ram[  673] = 'h000002a1; 	    data_ram[  674] = 'h000002a2; 	    data_ram[  675] = 'h000002a3; 	    data_ram[  676] = 'h000002a4; 	    data_ram[  677] = 'h000002a5; 	    data_ram[  678] = 'h000002a6; 	    data_ram[  679] = 'h000002a7; 	
    data_ram[  680] = 'h000002a8; 	    data_ram[  681] = 'h000002a9; 	    data_ram[  682] = 'h000002aa; 	    data_ram[  683] = 'h000002ab; 	    data_ram[  684] = 'h000002ac; 	    data_ram[  685] = 'h000002ad; 	    data_ram[  686] = 'h000002ae; 	    data_ram[  687] = 'h000002af; 	
    data_ram[  688] = 'h000002b0; 	    data_ram[  689] = 'h000002b1; 	    data_ram[  690] = 'h000002b2; 	    data_ram[  691] = 'h000002b3; 	    data_ram[  692] = 'h000002b4; 	    data_ram[  693] = 'h000002b5; 	    data_ram[  694] = 'h000002b6; 	    data_ram[  695] = 'h000002b7; 	
    data_ram[  696] = 'h000002b8; 	    data_ram[  697] = 'h000002b9; 	    data_ram[  698] = 'h000002ba; 	    data_ram[  699] = 'h000002bb; 	    data_ram[  700] = 'h000002bc; 	    data_ram[  701] = 'h000002bd; 	    data_ram[  702] = 'h000002be; 	    data_ram[  703] = 'h000002bf; 	
    data_ram[  704] = 'h000002c0; 	    data_ram[  705] = 'h000002c1; 	    data_ram[  706] = 'h000002c2; 	    data_ram[  707] = 'h000002c3; 	    data_ram[  708] = 'h000002c4; 	    data_ram[  709] = 'h000002c5; 	    data_ram[  710] = 'h000002c6; 	    data_ram[  711] = 'h000002c7; 	
    data_ram[  712] = 'h000002c8; 	    data_ram[  713] = 'h000002c9; 	    data_ram[  714] = 'h000002ca; 	    data_ram[  715] = 'h000002cb; 	    data_ram[  716] = 'h000002cc; 	    data_ram[  717] = 'h000002cd; 	    data_ram[  718] = 'h000002ce; 	    data_ram[  719] = 'h000002cf; 	
    data_ram[  720] = 'h000002d0; 	    data_ram[  721] = 'h000002d1; 	    data_ram[  722] = 'h000002d2; 	    data_ram[  723] = 'h000002d3; 	    data_ram[  724] = 'h000002d4; 	    data_ram[  725] = 'h000002d5; 	    data_ram[  726] = 'h000002d6; 	    data_ram[  727] = 'h000002d7; 	
    data_ram[  728] = 'h000002d8; 	    data_ram[  729] = 'h000002d9; 	    data_ram[  730] = 'h000002da; 	    data_ram[  731] = 'h000002db; 	    data_ram[  732] = 'h000002dc; 	    data_ram[  733] = 'h000002dd; 	    data_ram[  734] = 'h000002de; 	    data_ram[  735] = 'h000002df; 	
    data_ram[  736] = 'h000002e0; 	    data_ram[  737] = 'h000002e1; 	    data_ram[  738] = 'h000002e2; 	    data_ram[  739] = 'h000002e3; 	    data_ram[  740] = 'h000002e4; 	    data_ram[  741] = 'h000002e5; 	    data_ram[  742] = 'h000002e6; 	    data_ram[  743] = 'h000002e7; 	
    data_ram[  744] = 'h000002e8; 	    data_ram[  745] = 'h000002e9; 	    data_ram[  746] = 'h000002ea; 	    data_ram[  747] = 'h000002eb; 	    data_ram[  748] = 'h000002ec; 	    data_ram[  749] = 'h000002ed; 	    data_ram[  750] = 'h000002ee; 	    data_ram[  751] = 'h000002ef; 	
    data_ram[  752] = 'h000002f0; 	    data_ram[  753] = 'h000002f1; 	    data_ram[  754] = 'h000002f2; 	    data_ram[  755] = 'h000002f3; 	    data_ram[  756] = 'h000002f4; 	    data_ram[  757] = 'h000002f5; 	    data_ram[  758] = 'h000002f6; 	    data_ram[  759] = 'h000002f7; 	
    data_ram[  760] = 'h000002f8; 	    data_ram[  761] = 'h000002f9; 	    data_ram[  762] = 'h000002fa; 	    data_ram[  763] = 'h000002fb; 	    data_ram[  764] = 'h000002fc; 	    data_ram[  765] = 'h000002fd; 	    data_ram[  766] = 'h000002fe; 	    data_ram[  767] = 'h000002ff; 	
    data_ram[  768] = 'h00000300; 	    data_ram[  769] = 'h00000301; 	    data_ram[  770] = 'h00000302; 	    data_ram[  771] = 'h00000303; 	    data_ram[  772] = 'h00000304; 	    data_ram[  773] = 'h00000305; 	    data_ram[  774] = 'h00000306; 	    data_ram[  775] = 'h00000307; 	
    data_ram[  776] = 'h00000308; 	    data_ram[  777] = 'h00000309; 	    data_ram[  778] = 'h0000030a; 	    data_ram[  779] = 'h0000030b; 	    data_ram[  780] = 'h0000030c; 	    data_ram[  781] = 'h0000030d; 	    data_ram[  782] = 'h0000030e; 	    data_ram[  783] = 'h0000030f; 	
    data_ram[  784] = 'h00000310; 	    data_ram[  785] = 'h00000311; 	    data_ram[  786] = 'h00000312; 	    data_ram[  787] = 'h00000313; 	    data_ram[  788] = 'h00000314; 	    data_ram[  789] = 'h00000315; 	    data_ram[  790] = 'h00000316; 	    data_ram[  791] = 'h00000317; 	
    data_ram[  792] = 'h00000318; 	    data_ram[  793] = 'h00000319; 	    data_ram[  794] = 'h0000031a; 	    data_ram[  795] = 'h0000031b; 	    data_ram[  796] = 'h0000031c; 	    data_ram[  797] = 'h0000031d; 	    data_ram[  798] = 'h0000031e; 	    data_ram[  799] = 'h0000031f; 	
    data_ram[  800] = 'h00000320; 	    data_ram[  801] = 'h00000321; 	    data_ram[  802] = 'h00000322; 	    data_ram[  803] = 'h00000323; 	    data_ram[  804] = 'h00000324; 	    data_ram[  805] = 'h00000325; 	    data_ram[  806] = 'h00000326; 	    data_ram[  807] = 'h00000327; 	
    data_ram[  808] = 'h00000328; 	    data_ram[  809] = 'h00000329; 	    data_ram[  810] = 'h0000032a; 	    data_ram[  811] = 'h0000032b; 	    data_ram[  812] = 'h0000032c; 	    data_ram[  813] = 'h0000032d; 	    data_ram[  814] = 'h0000032e; 	    data_ram[  815] = 'h0000032f; 	
    data_ram[  816] = 'h00000330; 	    data_ram[  817] = 'h00000331; 	    data_ram[  818] = 'h00000332; 	    data_ram[  819] = 'h00000333; 	    data_ram[  820] = 'h00000334; 	    data_ram[  821] = 'h00000335; 	    data_ram[  822] = 'h00000336; 	    data_ram[  823] = 'h00000337; 	
    data_ram[  824] = 'h00000338; 	    data_ram[  825] = 'h00000339; 	    data_ram[  826] = 'h0000033a; 	    data_ram[  827] = 'h0000033b; 	    data_ram[  828] = 'h0000033c; 	    data_ram[  829] = 'h0000033d; 	    data_ram[  830] = 'h0000033e; 	    data_ram[  831] = 'h0000033f; 	
    data_ram[  832] = 'h00000340; 	    data_ram[  833] = 'h00000341; 	    data_ram[  834] = 'h00000342; 	    data_ram[  835] = 'h00000343; 	    data_ram[  836] = 'h00000344; 	    data_ram[  837] = 'h00000345; 	    data_ram[  838] = 'h00000346; 	    data_ram[  839] = 'h00000347; 	
    data_ram[  840] = 'h00000348; 	    data_ram[  841] = 'h00000349; 	    data_ram[  842] = 'h0000034a; 	    data_ram[  843] = 'h0000034b; 	    data_ram[  844] = 'h0000034c; 	    data_ram[  845] = 'h0000034d; 	    data_ram[  846] = 'h0000034e; 	    data_ram[  847] = 'h0000034f; 	
    data_ram[  848] = 'h00000350; 	    data_ram[  849] = 'h00000351; 	    data_ram[  850] = 'h00000352; 	    data_ram[  851] = 'h00000353; 	    data_ram[  852] = 'h00000354; 	    data_ram[  853] = 'h00000355; 	    data_ram[  854] = 'h00000356; 	    data_ram[  855] = 'h00000357; 	
    data_ram[  856] = 'h00000358; 	    data_ram[  857] = 'h00000359; 	    data_ram[  858] = 'h0000035a; 	    data_ram[  859] = 'h0000035b; 	    data_ram[  860] = 'h0000035c; 	    data_ram[  861] = 'h0000035d; 	    data_ram[  862] = 'h0000035e; 	    data_ram[  863] = 'h0000035f; 	
    data_ram[  864] = 'h00000360; 	    data_ram[  865] = 'h00000361; 	    data_ram[  866] = 'h00000362; 	    data_ram[  867] = 'h00000363; 	    data_ram[  868] = 'h00000364; 	    data_ram[  869] = 'h00000365; 	    data_ram[  870] = 'h00000366; 	    data_ram[  871] = 'h00000367; 	
    data_ram[  872] = 'h00000368; 	    data_ram[  873] = 'h00000369; 	    data_ram[  874] = 'h0000036a; 	    data_ram[  875] = 'h0000036b; 	    data_ram[  876] = 'h0000036c; 	    data_ram[  877] = 'h0000036d; 	    data_ram[  878] = 'h0000036e; 	    data_ram[  879] = 'h0000036f; 	
    data_ram[  880] = 'h00000370; 	    data_ram[  881] = 'h00000371; 	    data_ram[  882] = 'h00000372; 	    data_ram[  883] = 'h00000373; 	    data_ram[  884] = 'h00000374; 	    data_ram[  885] = 'h00000375; 	    data_ram[  886] = 'h00000376; 	    data_ram[  887] = 'h00000377; 	
    data_ram[  888] = 'h00000378; 	    data_ram[  889] = 'h00000379; 	    data_ram[  890] = 'h0000037a; 	    data_ram[  891] = 'h0000037b; 	    data_ram[  892] = 'h0000037c; 	    data_ram[  893] = 'h0000037d; 	    data_ram[  894] = 'h0000037e; 	    data_ram[  895] = 'h0000037f; 	
    data_ram[  896] = 'h00000380; 	    data_ram[  897] = 'h00000381; 	    data_ram[  898] = 'h00000382; 	    data_ram[  899] = 'h00000383; 	    data_ram[  900] = 'h00000384; 	    data_ram[  901] = 'h00000385; 	    data_ram[  902] = 'h00000386; 	    data_ram[  903] = 'h00000387; 	
    data_ram[  904] = 'h00000388; 	    data_ram[  905] = 'h00000389; 	    data_ram[  906] = 'h0000038a; 	    data_ram[  907] = 'h0000038b; 	    data_ram[  908] = 'h0000038c; 	    data_ram[  909] = 'h0000038d; 	    data_ram[  910] = 'h0000038e; 	    data_ram[  911] = 'h0000038f; 	
    data_ram[  912] = 'h00000390; 	    data_ram[  913] = 'h00000391; 	    data_ram[  914] = 'h00000392; 	    data_ram[  915] = 'h00000393; 	    data_ram[  916] = 'h00000394; 	    data_ram[  917] = 'h00000395; 	    data_ram[  918] = 'h00000396; 	    data_ram[  919] = 'h00000397; 	
    data_ram[  920] = 'h00000398; 	    data_ram[  921] = 'h00000399; 	    data_ram[  922] = 'h0000039a; 	    data_ram[  923] = 'h0000039b; 	    data_ram[  924] = 'h0000039c; 	    data_ram[  925] = 'h0000039d; 	    data_ram[  926] = 'h0000039e; 	    data_ram[  927] = 'h0000039f; 	
    data_ram[  928] = 'h000003a0; 	    data_ram[  929] = 'h000003a1; 	    data_ram[  930] = 'h000003a2; 	    data_ram[  931] = 'h000003a3; 	    data_ram[  932] = 'h000003a4; 	    data_ram[  933] = 'h000003a5; 	    data_ram[  934] = 'h000003a6; 	    data_ram[  935] = 'h000003a7; 	
    data_ram[  936] = 'h000003a8; 	    data_ram[  937] = 'h000003a9; 	    data_ram[  938] = 'h000003aa; 	    data_ram[  939] = 'h000003ab; 	    data_ram[  940] = 'h000003ac; 	    data_ram[  941] = 'h000003ad; 	    data_ram[  942] = 'h000003ae; 	    data_ram[  943] = 'h000003af; 	
    data_ram[  944] = 'h000003b0; 	    data_ram[  945] = 'h000003b1; 	    data_ram[  946] = 'h000003b2; 	    data_ram[  947] = 'h000003b3; 	    data_ram[  948] = 'h000003b4; 	    data_ram[  949] = 'h000003b5; 	    data_ram[  950] = 'h000003b6; 	    data_ram[  951] = 'h000003b7; 	
    data_ram[  952] = 'h000003b8; 	    data_ram[  953] = 'h000003b9; 	    data_ram[  954] = 'h000003ba; 	    data_ram[  955] = 'h000003bb; 	    data_ram[  956] = 'h000003bc; 	    data_ram[  957] = 'h000003bd; 	    data_ram[  958] = 'h000003be; 	    data_ram[  959] = 'h000003bf; 	
    data_ram[  960] = 'h000003c0; 	    data_ram[  961] = 'h000003c1; 	    data_ram[  962] = 'h000003c2; 	    data_ram[  963] = 'h000003c3; 	    data_ram[  964] = 'h000003c4; 	    data_ram[  965] = 'h000003c5; 	    data_ram[  966] = 'h000003c6; 	    data_ram[  967] = 'h000003c7; 	
    data_ram[  968] = 'h000003c8; 	    data_ram[  969] = 'h000003c9; 	    data_ram[  970] = 'h000003ca; 	    data_ram[  971] = 'h000003cb; 	    data_ram[  972] = 'h000003cc; 	    data_ram[  973] = 'h000003cd; 	    data_ram[  974] = 'h000003ce; 	    data_ram[  975] = 'h000003cf; 	
    data_ram[  976] = 'h000003d0; 	    data_ram[  977] = 'h000003d1; 	    data_ram[  978] = 'h000003d2; 	    data_ram[  979] = 'h000003d3; 	    data_ram[  980] = 'h000003d4; 	    data_ram[  981] = 'h000003d5; 	    data_ram[  982] = 'h000003d6; 	    data_ram[  983] = 'h000003d7; 	
    data_ram[  984] = 'h000003d8; 	    data_ram[  985] = 'h000003d9; 	    data_ram[  986] = 'h000003da; 	    data_ram[  987] = 'h000003db; 	    data_ram[  988] = 'h000003dc; 	    data_ram[  989] = 'h000003dd; 	    data_ram[  990] = 'h000003de; 	    data_ram[  991] = 'h000003df; 	
    data_ram[  992] = 'h000003e0; 	    data_ram[  993] = 'h000003e1; 	    data_ram[  994] = 'h000003e2; 	    data_ram[  995] = 'h000003e3; 	    data_ram[  996] = 'h000003e4; 	    data_ram[  997] = 'h000003e5; 	    data_ram[  998] = 'h000003e6; 	    data_ram[  999] = 'h000003e7; 	
    data_ram[ 1000] = 'h000003e8; 	    data_ram[ 1001] = 'h000003e9; 	    data_ram[ 1002] = 'h000003ea; 	    data_ram[ 1003] = 'h000003eb; 	    data_ram[ 1004] = 'h000003ec; 	    data_ram[ 1005] = 'h000003ed; 	    data_ram[ 1006] = 'h000003ee; 	    data_ram[ 1007] = 'h000003ef; 	
    data_ram[ 1008] = 'h000003f0; 	    data_ram[ 1009] = 'h000003f1; 	    data_ram[ 1010] = 'h000003f2; 	    data_ram[ 1011] = 'h000003f3; 	    data_ram[ 1012] = 'h000003f4; 	    data_ram[ 1013] = 'h000003f5; 	    data_ram[ 1014] = 'h000003f6; 	    data_ram[ 1015] = 'h000003f7; 	
    data_ram[ 1016] = 'h000003f8; 	    data_ram[ 1017] = 'h000003f9; 	    data_ram[ 1018] = 'h000003fa; 	    data_ram[ 1019] = 'h000003fb; 	    data_ram[ 1020] = 'h000003fc; 	    data_ram[ 1021] = 'h000003fd; 	    data_ram[ 1022] = 'h000003fe; 	    data_ram[ 1023] = 'h000003ff; 	

end
initial begin
    i_addr_rom[    0] = 'h0000009c; 	    d_addr_rom[    0] = 'h000008b8; 	    wdata_rom[    0] = 'h53936e4e; 	    wvalid_rom[    0] = 0; 
    i_addr_rom[    1] = 'h00000540; 	    d_addr_rom[    1] = 'h0000094c; 	    wdata_rom[    1] = 'h152428b1; 	    wvalid_rom[    1] = 1; 
    i_addr_rom[    2] = 'h000003fc; 	    d_addr_rom[    2] = 'h00000d08; 	    wdata_rom[    2] = 'heb6d07be; 	    wvalid_rom[    2] = 0; 
    i_addr_rom[    3] = 'h00000118; 	    d_addr_rom[    3] = 'h0000085c; 	    wdata_rom[    3] = 'hb01f3cb4; 	    wvalid_rom[    3] = 1; 
    i_addr_rom[    4] = 'h000000e4; 	    d_addr_rom[    4] = 'h00000e10; 	    wdata_rom[    4] = 'hcc0f0c59; 	    wvalid_rom[    4] = 0; 
    i_addr_rom[    5] = 'h00000290; 	    d_addr_rom[    5] = 'h00000bdc; 	    wdata_rom[    5] = 'h95ca3206; 	    wvalid_rom[    5] = 0; 
    i_addr_rom[    6] = 'h000001a8; 	    d_addr_rom[    6] = 'h00000d8c; 	    wdata_rom[    6] = 'ha116ab10; 	    wvalid_rom[    6] = 1; 
    i_addr_rom[    7] = 'h00000758; 	    d_addr_rom[    7] = 'h00000dbc; 	    wdata_rom[    7] = 'h6a70cd11; 	    wvalid_rom[    7] = 0; 
    i_addr_rom[    8] = 'h00000424; 	    d_addr_rom[    8] = 'h00000d44; 	    wdata_rom[    8] = 'h9c098e68; 	    wvalid_rom[    8] = 1; 
    i_addr_rom[    9] = 'h000000a8; 	    d_addr_rom[    9] = 'h00000e6c; 	    wdata_rom[    9] = 'h2a51bcb6; 	    wvalid_rom[    9] = 1; 
    i_addr_rom[   10] = 'h00000218; 	    d_addr_rom[   10] = 'h00000c08; 	    wdata_rom[   10] = 'h6c241477; 	    wvalid_rom[   10] = 0; 
    i_addr_rom[   11] = 'h00000730; 	    d_addr_rom[   11] = 'h00000bdc; 	    wdata_rom[   11] = 'h9eb6e356; 	    wvalid_rom[   11] = 1; 
    i_addr_rom[   12] = 'h0000019c; 	    d_addr_rom[   12] = 'h00000ba8; 	    wdata_rom[   12] = 'h180e298d; 	    wvalid_rom[   12] = 1; 
    i_addr_rom[   13] = 'h000001f0; 	    d_addr_rom[   13] = 'h00000dc4; 	    wdata_rom[   13] = 'h0140d5d0; 	    wvalid_rom[   13] = 1; 
    i_addr_rom[   14] = 'h00000278; 	    d_addr_rom[   14] = 'h00000874; 	    wdata_rom[   14] = 'h23b071f3; 	    wvalid_rom[   14] = 1; 
    i_addr_rom[   15] = 'h00000778; 	    d_addr_rom[   15] = 'h000009e0; 	    wdata_rom[   15] = 'h68fb60c1; 	    wvalid_rom[   15] = 0; 
    i_addr_rom[   16] = 'h00000394; 	    d_addr_rom[   16] = 'h000009b0; 	    wdata_rom[   16] = 'h4f317ae4; 	    wvalid_rom[   16] = 1; 
    i_addr_rom[   17] = 'h0000079c; 	    d_addr_rom[   17] = 'h00000ec0; 	    wdata_rom[   17] = 'hb2d356fe; 	    wvalid_rom[   17] = 1; 
    i_addr_rom[   18] = 'h000000f0; 	    d_addr_rom[   18] = 'h00000a20; 	    wdata_rom[   18] = 'h99971305; 	    wvalid_rom[   18] = 1; 
    i_addr_rom[   19] = 'h000001d0; 	    d_addr_rom[   19] = 'h000009c8; 	    wdata_rom[   19] = 'haffa59a1; 	    wvalid_rom[   19] = 1; 
    i_addr_rom[   20] = 'h000001a4; 	    d_addr_rom[   20] = 'h000009d8; 	    wdata_rom[   20] = 'h7a520bba; 	    wvalid_rom[   20] = 1; 
    i_addr_rom[   21] = 'h0000076c; 	    d_addr_rom[   21] = 'h00000b34; 	    wdata_rom[   21] = 'h67f5b96a; 	    wvalid_rom[   21] = 0; 
    i_addr_rom[   22] = 'h00000178; 	    d_addr_rom[   22] = 'h00000aa4; 	    wdata_rom[   22] = 'h0f64aa62; 	    wvalid_rom[   22] = 1; 
    i_addr_rom[   23] = 'h00000204; 	    d_addr_rom[   23] = 'h00000d28; 	    wdata_rom[   23] = 'hb02eb24a; 	    wvalid_rom[   23] = 0; 
    i_addr_rom[   24] = 'h00000448; 	    d_addr_rom[   24] = 'h00000a6c; 	    wdata_rom[   24] = 'h07b821f6; 	    wvalid_rom[   24] = 1; 
    i_addr_rom[   25] = 'h0000046c; 	    d_addr_rom[   25] = 'h00000f34; 	    wdata_rom[   25] = 'h0aad9093; 	    wvalid_rom[   25] = 1; 
    i_addr_rom[   26] = 'h00000204; 	    d_addr_rom[   26] = 'h00000db4; 	    wdata_rom[   26] = 'h72f94911; 	    wvalid_rom[   26] = 1; 
    i_addr_rom[   27] = 'h00000350; 	    d_addr_rom[   27] = 'h00000f50; 	    wdata_rom[   27] = 'h5b1ef34f; 	    wvalid_rom[   27] = 1; 
    i_addr_rom[   28] = 'h00000028; 	    d_addr_rom[   28] = 'h00000c98; 	    wdata_rom[   28] = 'hf12f5240; 	    wvalid_rom[   28] = 0; 
    i_addr_rom[   29] = 'h000006e4; 	    d_addr_rom[   29] = 'h00000cc8; 	    wdata_rom[   29] = 'h92a51691; 	    wvalid_rom[   29] = 1; 
    i_addr_rom[   30] = 'h00000504; 	    d_addr_rom[   30] = 'h00000ff0; 	    wdata_rom[   30] = 'hf3f84584; 	    wvalid_rom[   30] = 0; 
    i_addr_rom[   31] = 'h000003c8; 	    d_addr_rom[   31] = 'h00000adc; 	    wdata_rom[   31] = 'h424a299b; 	    wvalid_rom[   31] = 1; 
    i_addr_rom[   32] = 'h0000047c; 	    d_addr_rom[   32] = 'h00000e00; 	    wdata_rom[   32] = 'h3b51669b; 	    wvalid_rom[   32] = 0; 
    i_addr_rom[   33] = 'h00000510; 	    d_addr_rom[   33] = 'h00000cc0; 	    wdata_rom[   33] = 'h34c44d29; 	    wvalid_rom[   33] = 1; 
    i_addr_rom[   34] = 'h0000007c; 	    d_addr_rom[   34] = 'h00000e08; 	    wdata_rom[   34] = 'ha2fdf764; 	    wvalid_rom[   34] = 0; 
    i_addr_rom[   35] = 'h00000644; 	    d_addr_rom[   35] = 'h00000a20; 	    wdata_rom[   35] = 'ha1b1474f; 	    wvalid_rom[   35] = 0; 
    i_addr_rom[   36] = 'h000007f8; 	    d_addr_rom[   36] = 'h00000ca0; 	    wdata_rom[   36] = 'h3870b079; 	    wvalid_rom[   36] = 0; 
    i_addr_rom[   37] = 'h00000218; 	    d_addr_rom[   37] = 'h00000840; 	    wdata_rom[   37] = 'h82ab6bf0; 	    wvalid_rom[   37] = 1; 
    i_addr_rom[   38] = 'h00000290; 	    d_addr_rom[   38] = 'h00000adc; 	    wdata_rom[   38] = 'h9ba50c16; 	    wvalid_rom[   38] = 1; 
    i_addr_rom[   39] = 'h0000025c; 	    d_addr_rom[   39] = 'h00000b2c; 	    wdata_rom[   39] = 'h58d10490; 	    wvalid_rom[   39] = 1; 
    i_addr_rom[   40] = 'h000003bc; 	    d_addr_rom[   40] = 'h00000f48; 	    wdata_rom[   40] = 'h40f582ad; 	    wvalid_rom[   40] = 1; 
    i_addr_rom[   41] = 'h000000fc; 	    d_addr_rom[   41] = 'h000008b0; 	    wdata_rom[   41] = 'h6cff2b55; 	    wvalid_rom[   41] = 0; 
    i_addr_rom[   42] = 'h000005cc; 	    d_addr_rom[   42] = 'h00000db8; 	    wdata_rom[   42] = 'h9ba6a68e; 	    wvalid_rom[   42] = 0; 
    i_addr_rom[   43] = 'h0000023c; 	    d_addr_rom[   43] = 'h00000f80; 	    wdata_rom[   43] = 'ha9fbf25b; 	    wvalid_rom[   43] = 0; 
    i_addr_rom[   44] = 'h000005e4; 	    d_addr_rom[   44] = 'h000008b8; 	    wdata_rom[   44] = 'h60f6df94; 	    wvalid_rom[   44] = 0; 
    i_addr_rom[   45] = 'h00000434; 	    d_addr_rom[   45] = 'h00000e04; 	    wdata_rom[   45] = 'h0314c48f; 	    wvalid_rom[   45] = 1; 
    i_addr_rom[   46] = 'h00000444; 	    d_addr_rom[   46] = 'h000009c4; 	    wdata_rom[   46] = 'h3543fcc9; 	    wvalid_rom[   46] = 0; 
    i_addr_rom[   47] = 'h000004e0; 	    d_addr_rom[   47] = 'h00000cfc; 	    wdata_rom[   47] = 'hbee6ac52; 	    wvalid_rom[   47] = 1; 
    i_addr_rom[   48] = 'h0000035c; 	    d_addr_rom[   48] = 'h00000a68; 	    wdata_rom[   48] = 'hb710cf32; 	    wvalid_rom[   48] = 0; 
    i_addr_rom[   49] = 'h000005c0; 	    d_addr_rom[   49] = 'h00000b64; 	    wdata_rom[   49] = 'h9ef3b268; 	    wvalid_rom[   49] = 0; 
    i_addr_rom[   50] = 'h000000e8; 	    d_addr_rom[   50] = 'h00000c04; 	    wdata_rom[   50] = 'h355a4ff7; 	    wvalid_rom[   50] = 0; 
    i_addr_rom[   51] = 'h000005a4; 	    d_addr_rom[   51] = 'h00000a78; 	    wdata_rom[   51] = 'h5d1746c4; 	    wvalid_rom[   51] = 1; 
    i_addr_rom[   52] = 'h000000a8; 	    d_addr_rom[   52] = 'h000008a0; 	    wdata_rom[   52] = 'h6ebb5d1c; 	    wvalid_rom[   52] = 1; 
    i_addr_rom[   53] = 'h00000400; 	    d_addr_rom[   53] = 'h00000fb4; 	    wdata_rom[   53] = 'hc77ab386; 	    wvalid_rom[   53] = 0; 
    i_addr_rom[   54] = 'h000000b8; 	    d_addr_rom[   54] = 'h00000d88; 	    wdata_rom[   54] = 'h05755dcb; 	    wvalid_rom[   54] = 1; 
    i_addr_rom[   55] = 'h00000720; 	    d_addr_rom[   55] = 'h00000bf0; 	    wdata_rom[   55] = 'h9b45a1c8; 	    wvalid_rom[   55] = 0; 
    i_addr_rom[   56] = 'h000002e0; 	    d_addr_rom[   56] = 'h00000fb8; 	    wdata_rom[   56] = 'h58b69500; 	    wvalid_rom[   56] = 0; 
    i_addr_rom[   57] = 'h00000088; 	    d_addr_rom[   57] = 'h0000090c; 	    wdata_rom[   57] = 'hd43c94a6; 	    wvalid_rom[   57] = 1; 
    i_addr_rom[   58] = 'h000006ec; 	    d_addr_rom[   58] = 'h00000e3c; 	    wdata_rom[   58] = 'h68d170d0; 	    wvalid_rom[   58] = 1; 
    i_addr_rom[   59] = 'h00000264; 	    d_addr_rom[   59] = 'h00000aa0; 	    wdata_rom[   59] = 'hb4dd2d66; 	    wvalid_rom[   59] = 0; 
    i_addr_rom[   60] = 'h000005f8; 	    d_addr_rom[   60] = 'h00000ac4; 	    wdata_rom[   60] = 'h3263ec05; 	    wvalid_rom[   60] = 0; 
    i_addr_rom[   61] = 'h00000594; 	    d_addr_rom[   61] = 'h00000cc4; 	    wdata_rom[   61] = 'hc636116b; 	    wvalid_rom[   61] = 0; 
    i_addr_rom[   62] = 'h000003ec; 	    d_addr_rom[   62] = 'h000009d0; 	    wdata_rom[   62] = 'h6baf133b; 	    wvalid_rom[   62] = 1; 
    i_addr_rom[   63] = 'h00000764; 	    d_addr_rom[   63] = 'h00000da8; 	    wdata_rom[   63] = 'hf9542bbc; 	    wvalid_rom[   63] = 0; 
    i_addr_rom[   64] = 'h000006d8; 	    d_addr_rom[   64] = 'h00000a94; 	    wdata_rom[   64] = 'h4c769b7f; 	    wvalid_rom[   64] = 1; 
    i_addr_rom[   65] = 'h000006dc; 	    d_addr_rom[   65] = 'h00000c30; 	    wdata_rom[   65] = 'h60a11cc1; 	    wvalid_rom[   65] = 0; 
    i_addr_rom[   66] = 'h00000790; 	    d_addr_rom[   66] = 'h00000c30; 	    wdata_rom[   66] = 'h0e72051a; 	    wvalid_rom[   66] = 1; 
    i_addr_rom[   67] = 'h000005d8; 	    d_addr_rom[   67] = 'h000009c4; 	    wdata_rom[   67] = 'h492d51d0; 	    wvalid_rom[   67] = 0; 
    i_addr_rom[   68] = 'h00000334; 	    d_addr_rom[   68] = 'h00000b08; 	    wdata_rom[   68] = 'h68225c1b; 	    wvalid_rom[   68] = 1; 
    i_addr_rom[   69] = 'h000005fc; 	    d_addr_rom[   69] = 'h00000ca0; 	    wdata_rom[   69] = 'hc10cf127; 	    wvalid_rom[   69] = 1; 
    i_addr_rom[   70] = 'h000000b0; 	    d_addr_rom[   70] = 'h000008cc; 	    wdata_rom[   70] = 'h306a96f0; 	    wvalid_rom[   70] = 1; 
    i_addr_rom[   71] = 'h000001d4; 	    d_addr_rom[   71] = 'h00000858; 	    wdata_rom[   71] = 'h89c5cb1d; 	    wvalid_rom[   71] = 0; 
    i_addr_rom[   72] = 'h00000024; 	    d_addr_rom[   72] = 'h00000ac8; 	    wdata_rom[   72] = 'h534f6612; 	    wvalid_rom[   72] = 0; 
    i_addr_rom[   73] = 'h000007b8; 	    d_addr_rom[   73] = 'h00000fe8; 	    wdata_rom[   73] = 'h659425b8; 	    wvalid_rom[   73] = 0; 
    i_addr_rom[   74] = 'h0000016c; 	    d_addr_rom[   74] = 'h00000b94; 	    wdata_rom[   74] = 'hcb086723; 	    wvalid_rom[   74] = 1; 
    i_addr_rom[   75] = 'h000006f0; 	    d_addr_rom[   75] = 'h00000b6c; 	    wdata_rom[   75] = 'h20a30a22; 	    wvalid_rom[   75] = 1; 
    i_addr_rom[   76] = 'h00000508; 	    d_addr_rom[   76] = 'h00000f80; 	    wdata_rom[   76] = 'h8c1c8d6e; 	    wvalid_rom[   76] = 0; 
    i_addr_rom[   77] = 'h000007e4; 	    d_addr_rom[   77] = 'h00000ef4; 	    wdata_rom[   77] = 'h3e5a8021; 	    wvalid_rom[   77] = 0; 
    i_addr_rom[   78] = 'h000007e0; 	    d_addr_rom[   78] = 'h00000f10; 	    wdata_rom[   78] = 'h769d68c1; 	    wvalid_rom[   78] = 0; 
    i_addr_rom[   79] = 'h000000a0; 	    d_addr_rom[   79] = 'h00000d98; 	    wdata_rom[   79] = 'h08829a02; 	    wvalid_rom[   79] = 1; 
    i_addr_rom[   80] = 'h000005f8; 	    d_addr_rom[   80] = 'h00000da0; 	    wdata_rom[   80] = 'h0a08a4bf; 	    wvalid_rom[   80] = 0; 
    i_addr_rom[   81] = 'h00000128; 	    d_addr_rom[   81] = 'h00000efc; 	    wdata_rom[   81] = 'hbe3d9387; 	    wvalid_rom[   81] = 0; 
    i_addr_rom[   82] = 'h000004e0; 	    d_addr_rom[   82] = 'h00000c04; 	    wdata_rom[   82] = 'hb0fc362c; 	    wvalid_rom[   82] = 0; 
    i_addr_rom[   83] = 'h000006c4; 	    d_addr_rom[   83] = 'h00000b68; 	    wdata_rom[   83] = 'h0903bd26; 	    wvalid_rom[   83] = 1; 
    i_addr_rom[   84] = 'h000000d0; 	    d_addr_rom[   84] = 'h00000c78; 	    wdata_rom[   84] = 'h3b6c3383; 	    wvalid_rom[   84] = 0; 
    i_addr_rom[   85] = 'h000005f0; 	    d_addr_rom[   85] = 'h000009d0; 	    wdata_rom[   85] = 'h52ae796f; 	    wvalid_rom[   85] = 1; 
    i_addr_rom[   86] = 'h00000684; 	    d_addr_rom[   86] = 'h00000b28; 	    wdata_rom[   86] = 'hdd2aef25; 	    wvalid_rom[   86] = 1; 
    i_addr_rom[   87] = 'h00000378; 	    d_addr_rom[   87] = 'h00000834; 	    wdata_rom[   87] = 'h2a9817cc; 	    wvalid_rom[   87] = 0; 
    i_addr_rom[   88] = 'h00000008; 	    d_addr_rom[   88] = 'h00000e3c; 	    wdata_rom[   88] = 'h804fb81a; 	    wvalid_rom[   88] = 0; 
    i_addr_rom[   89] = 'h0000025c; 	    d_addr_rom[   89] = 'h00000b48; 	    wdata_rom[   89] = 'h96a158a5; 	    wvalid_rom[   89] = 1; 
    i_addr_rom[   90] = 'h00000314; 	    d_addr_rom[   90] = 'h00000d64; 	    wdata_rom[   90] = 'hfb1b3733; 	    wvalid_rom[   90] = 1; 
    i_addr_rom[   91] = 'h00000068; 	    d_addr_rom[   91] = 'h00000a00; 	    wdata_rom[   91] = 'ha6c2e57c; 	    wvalid_rom[   91] = 0; 
    i_addr_rom[   92] = 'h00000294; 	    d_addr_rom[   92] = 'h00000ccc; 	    wdata_rom[   92] = 'h2100b8c6; 	    wvalid_rom[   92] = 0; 
    i_addr_rom[   93] = 'h00000784; 	    d_addr_rom[   93] = 'h00000c10; 	    wdata_rom[   93] = 'hf3931991; 	    wvalid_rom[   93] = 1; 
    i_addr_rom[   94] = 'h0000075c; 	    d_addr_rom[   94] = 'h00000e88; 	    wdata_rom[   94] = 'h419f1d84; 	    wvalid_rom[   94] = 0; 
    i_addr_rom[   95] = 'h00000524; 	    d_addr_rom[   95] = 'h00000bbc; 	    wdata_rom[   95] = 'hacdae3a3; 	    wvalid_rom[   95] = 1; 
    i_addr_rom[   96] = 'h00000074; 	    d_addr_rom[   96] = 'h00000f60; 	    wdata_rom[   96] = 'ha8e0600b; 	    wvalid_rom[   96] = 0; 
    i_addr_rom[   97] = 'h000004b0; 	    d_addr_rom[   97] = 'h00000ee0; 	    wdata_rom[   97] = 'h6a9514ad; 	    wvalid_rom[   97] = 0; 
    i_addr_rom[   98] = 'h00000574; 	    d_addr_rom[   98] = 'h00000dc4; 	    wdata_rom[   98] = 'hb5997cc8; 	    wvalid_rom[   98] = 0; 
    i_addr_rom[   99] = 'h00000734; 	    d_addr_rom[   99] = 'h00000a28; 	    wdata_rom[   99] = 'h705708c9; 	    wvalid_rom[   99] = 1; 
    i_addr_rom[  100] = 'h00000044; 	    d_addr_rom[  100] = 'h00000c20; 	    wdata_rom[  100] = 'h10803dff; 	    wvalid_rom[  100] = 0; 
    i_addr_rom[  101] = 'h00000070; 	    d_addr_rom[  101] = 'h00000d64; 	    wdata_rom[  101] = 'hdca64147; 	    wvalid_rom[  101] = 0; 
    i_addr_rom[  102] = 'h00000040; 	    d_addr_rom[  102] = 'h0000087c; 	    wdata_rom[  102] = 'h3505a3ed; 	    wvalid_rom[  102] = 1; 
    i_addr_rom[  103] = 'h000003b4; 	    d_addr_rom[  103] = 'h000009a0; 	    wdata_rom[  103] = 'hb40e7ca3; 	    wvalid_rom[  103] = 1; 
    i_addr_rom[  104] = 'h000001dc; 	    d_addr_rom[  104] = 'h00000b04; 	    wdata_rom[  104] = 'h07484bf7; 	    wvalid_rom[  104] = 1; 
    i_addr_rom[  105] = 'h00000730; 	    d_addr_rom[  105] = 'h00000af8; 	    wdata_rom[  105] = 'hb64133bb; 	    wvalid_rom[  105] = 0; 
    i_addr_rom[  106] = 'h0000037c; 	    d_addr_rom[  106] = 'h00000904; 	    wdata_rom[  106] = 'h65a48908; 	    wvalid_rom[  106] = 1; 
    i_addr_rom[  107] = 'h0000020c; 	    d_addr_rom[  107] = 'h00000c3c; 	    wdata_rom[  107] = 'h7cd0d098; 	    wvalid_rom[  107] = 1; 
    i_addr_rom[  108] = 'h00000660; 	    d_addr_rom[  108] = 'h00000878; 	    wdata_rom[  108] = 'h7da4a53e; 	    wvalid_rom[  108] = 1; 
    i_addr_rom[  109] = 'h0000008c; 	    d_addr_rom[  109] = 'h00000d78; 	    wdata_rom[  109] = 'hbe62b07f; 	    wvalid_rom[  109] = 0; 
    i_addr_rom[  110] = 'h00000418; 	    d_addr_rom[  110] = 'h00000b00; 	    wdata_rom[  110] = 'h859b2656; 	    wvalid_rom[  110] = 0; 
    i_addr_rom[  111] = 'h000000c4; 	    d_addr_rom[  111] = 'h00000c34; 	    wdata_rom[  111] = 'h970e8080; 	    wvalid_rom[  111] = 0; 
    i_addr_rom[  112] = 'h000004f4; 	    d_addr_rom[  112] = 'h00000ea4; 	    wdata_rom[  112] = 'hd52aad5f; 	    wvalid_rom[  112] = 0; 
    i_addr_rom[  113] = 'h000006f0; 	    d_addr_rom[  113] = 'h00000a70; 	    wdata_rom[  113] = 'hbb94a81b; 	    wvalid_rom[  113] = 0; 
    i_addr_rom[  114] = 'h000002d0; 	    d_addr_rom[  114] = 'h00000df8; 	    wdata_rom[  114] = 'h847e1fb3; 	    wvalid_rom[  114] = 0; 
    i_addr_rom[  115] = 'h00000378; 	    d_addr_rom[  115] = 'h00000dc0; 	    wdata_rom[  115] = 'h70e3d755; 	    wvalid_rom[  115] = 1; 
    i_addr_rom[  116] = 'h00000744; 	    d_addr_rom[  116] = 'h00000d14; 	    wdata_rom[  116] = 'h238d711d; 	    wvalid_rom[  116] = 0; 
    i_addr_rom[  117] = 'h0000056c; 	    d_addr_rom[  117] = 'h00000a7c; 	    wdata_rom[  117] = 'h61b86c75; 	    wvalid_rom[  117] = 0; 
    i_addr_rom[  118] = 'h000000a8; 	    d_addr_rom[  118] = 'h0000091c; 	    wdata_rom[  118] = 'h224dd823; 	    wvalid_rom[  118] = 0; 
    i_addr_rom[  119] = 'h00000288; 	    d_addr_rom[  119] = 'h00000f00; 	    wdata_rom[  119] = 'hff64cd24; 	    wvalid_rom[  119] = 1; 
    i_addr_rom[  120] = 'h00000194; 	    d_addr_rom[  120] = 'h00000924; 	    wdata_rom[  120] = 'he4d873a4; 	    wvalid_rom[  120] = 1; 
    i_addr_rom[  121] = 'h0000064c; 	    d_addr_rom[  121] = 'h00000c88; 	    wdata_rom[  121] = 'h001ae3ca; 	    wvalid_rom[  121] = 1; 
    i_addr_rom[  122] = 'h000002a0; 	    d_addr_rom[  122] = 'h00000a98; 	    wdata_rom[  122] = 'ha8a81d18; 	    wvalid_rom[  122] = 1; 
    i_addr_rom[  123] = 'h000000e8; 	    d_addr_rom[  123] = 'h00000840; 	    wdata_rom[  123] = 'h022dc689; 	    wvalid_rom[  123] = 0; 
    i_addr_rom[  124] = 'h000007f0; 	    d_addr_rom[  124] = 'h00000a24; 	    wdata_rom[  124] = 'hff93847c; 	    wvalid_rom[  124] = 0; 
    i_addr_rom[  125] = 'h0000011c; 	    d_addr_rom[  125] = 'h00000f00; 	    wdata_rom[  125] = 'h5f8501f6; 	    wvalid_rom[  125] = 1; 
    i_addr_rom[  126] = 'h00000250; 	    d_addr_rom[  126] = 'h00000930; 	    wdata_rom[  126] = 'h1fd88b97; 	    wvalid_rom[  126] = 1; 
    i_addr_rom[  127] = 'h000003e4; 	    d_addr_rom[  127] = 'h00000cfc; 	    wdata_rom[  127] = 'hb51dbbb8; 	    wvalid_rom[  127] = 1; 
    i_addr_rom[  128] = 'h00000488; 	    d_addr_rom[  128] = 'h00000d94; 	    wdata_rom[  128] = 'h2f2347cd; 	    wvalid_rom[  128] = 0; 
    i_addr_rom[  129] = 'h000002f4; 	    d_addr_rom[  129] = 'h000009e8; 	    wdata_rom[  129] = 'h1a45d974; 	    wvalid_rom[  129] = 0; 
    i_addr_rom[  130] = 'h000007a4; 	    d_addr_rom[  130] = 'h00000c04; 	    wdata_rom[  130] = 'hf2fad0fa; 	    wvalid_rom[  130] = 0; 
    i_addr_rom[  131] = 'h00000724; 	    d_addr_rom[  131] = 'h00000a30; 	    wdata_rom[  131] = 'hc05d0b39; 	    wvalid_rom[  131] = 0; 
    i_addr_rom[  132] = 'h00000700; 	    d_addr_rom[  132] = 'h00000df4; 	    wdata_rom[  132] = 'ha2703b2e; 	    wvalid_rom[  132] = 0; 
    i_addr_rom[  133] = 'h000004d8; 	    d_addr_rom[  133] = 'h00000ea4; 	    wdata_rom[  133] = 'hffeb0900; 	    wvalid_rom[  133] = 1; 
    i_addr_rom[  134] = 'h000003cc; 	    d_addr_rom[  134] = 'h00000c9c; 	    wdata_rom[  134] = 'h2b156884; 	    wvalid_rom[  134] = 1; 
    i_addr_rom[  135] = 'h00000708; 	    d_addr_rom[  135] = 'h00000958; 	    wdata_rom[  135] = 'hd710da75; 	    wvalid_rom[  135] = 1; 
    i_addr_rom[  136] = 'h0000010c; 	    d_addr_rom[  136] = 'h00000c7c; 	    wdata_rom[  136] = 'hc77cefef; 	    wvalid_rom[  136] = 0; 
    i_addr_rom[  137] = 'h0000044c; 	    d_addr_rom[  137] = 'h00000c44; 	    wdata_rom[  137] = 'ha08924ec; 	    wvalid_rom[  137] = 1; 
    i_addr_rom[  138] = 'h0000020c; 	    d_addr_rom[  138] = 'h00000a9c; 	    wdata_rom[  138] = 'he92f6131; 	    wvalid_rom[  138] = 0; 
    i_addr_rom[  139] = 'h00000604; 	    d_addr_rom[  139] = 'h00000ef4; 	    wdata_rom[  139] = 'hddc2f82a; 	    wvalid_rom[  139] = 0; 
    i_addr_rom[  140] = 'h00000468; 	    d_addr_rom[  140] = 'h00000cac; 	    wdata_rom[  140] = 'h955e60f2; 	    wvalid_rom[  140] = 0; 
    i_addr_rom[  141] = 'h00000404; 	    d_addr_rom[  141] = 'h00000958; 	    wdata_rom[  141] = 'h34e4221d; 	    wvalid_rom[  141] = 0; 
    i_addr_rom[  142] = 'h000002ec; 	    d_addr_rom[  142] = 'h00000eb8; 	    wdata_rom[  142] = 'hd0f86e7f; 	    wvalid_rom[  142] = 1; 
    i_addr_rom[  143] = 'h000000d4; 	    d_addr_rom[  143] = 'h00000a10; 	    wdata_rom[  143] = 'h02d767d4; 	    wvalid_rom[  143] = 1; 
    i_addr_rom[  144] = 'h00000728; 	    d_addr_rom[  144] = 'h00000b08; 	    wdata_rom[  144] = 'hd6164c18; 	    wvalid_rom[  144] = 0; 
    i_addr_rom[  145] = 'h000000fc; 	    d_addr_rom[  145] = 'h00000894; 	    wdata_rom[  145] = 'h875b6527; 	    wvalid_rom[  145] = 0; 
    i_addr_rom[  146] = 'h00000730; 	    d_addr_rom[  146] = 'h00000de4; 	    wdata_rom[  146] = 'h619a26b1; 	    wvalid_rom[  146] = 1; 
    i_addr_rom[  147] = 'h0000076c; 	    d_addr_rom[  147] = 'h00000d64; 	    wdata_rom[  147] = 'h62230ccb; 	    wvalid_rom[  147] = 1; 
    i_addr_rom[  148] = 'h000002ec; 	    d_addr_rom[  148] = 'h00000e34; 	    wdata_rom[  148] = 'h42c8e97d; 	    wvalid_rom[  148] = 0; 
    i_addr_rom[  149] = 'h00000430; 	    d_addr_rom[  149] = 'h00000e58; 	    wdata_rom[  149] = 'h2c7e3e03; 	    wvalid_rom[  149] = 0; 
    i_addr_rom[  150] = 'h00000474; 	    d_addr_rom[  150] = 'h00000bac; 	    wdata_rom[  150] = 'hedf79ab7; 	    wvalid_rom[  150] = 0; 
    i_addr_rom[  151] = 'h000005ac; 	    d_addr_rom[  151] = 'h00000fdc; 	    wdata_rom[  151] = 'h63d171be; 	    wvalid_rom[  151] = 1; 
    i_addr_rom[  152] = 'h000005cc; 	    d_addr_rom[  152] = 'h00000990; 	    wdata_rom[  152] = 'h769491eb; 	    wvalid_rom[  152] = 1; 
    i_addr_rom[  153] = 'h00000218; 	    d_addr_rom[  153] = 'h00000ba8; 	    wdata_rom[  153] = 'h21328c8d; 	    wvalid_rom[  153] = 0; 
    i_addr_rom[  154] = 'h00000738; 	    d_addr_rom[  154] = 'h00000804; 	    wdata_rom[  154] = 'h7cf7abf8; 	    wvalid_rom[  154] = 0; 
    i_addr_rom[  155] = 'h000002b4; 	    d_addr_rom[  155] = 'h00000818; 	    wdata_rom[  155] = 'hfeb900bd; 	    wvalid_rom[  155] = 0; 
    i_addr_rom[  156] = 'h00000620; 	    d_addr_rom[  156] = 'h00000fc8; 	    wdata_rom[  156] = 'hc12002d5; 	    wvalid_rom[  156] = 0; 
    i_addr_rom[  157] = 'h000002ac; 	    d_addr_rom[  157] = 'h00000848; 	    wdata_rom[  157] = 'h7bb446df; 	    wvalid_rom[  157] = 0; 
    i_addr_rom[  158] = 'h000006ac; 	    d_addr_rom[  158] = 'h00000fe8; 	    wdata_rom[  158] = 'h749d7bb0; 	    wvalid_rom[  158] = 0; 
    i_addr_rom[  159] = 'h0000004c; 	    d_addr_rom[  159] = 'h00000da0; 	    wdata_rom[  159] = 'hdee3c705; 	    wvalid_rom[  159] = 1; 
    i_addr_rom[  160] = 'h000003a0; 	    d_addr_rom[  160] = 'h00000e98; 	    wdata_rom[  160] = 'h1cdc56e8; 	    wvalid_rom[  160] = 1; 
    i_addr_rom[  161] = 'h000006c4; 	    d_addr_rom[  161] = 'h00000f38; 	    wdata_rom[  161] = 'hc3e20a61; 	    wvalid_rom[  161] = 1; 
    i_addr_rom[  162] = 'h00000050; 	    d_addr_rom[  162] = 'h00000bf4; 	    wdata_rom[  162] = 'h0c64cf51; 	    wvalid_rom[  162] = 0; 
    i_addr_rom[  163] = 'h0000044c; 	    d_addr_rom[  163] = 'h00000c60; 	    wdata_rom[  163] = 'h17481d66; 	    wvalid_rom[  163] = 1; 
    i_addr_rom[  164] = 'h000000f4; 	    d_addr_rom[  164] = 'h00000fdc; 	    wdata_rom[  164] = 'he20b4ef0; 	    wvalid_rom[  164] = 1; 
    i_addr_rom[  165] = 'h00000160; 	    d_addr_rom[  165] = 'h00000eec; 	    wdata_rom[  165] = 'hdaf144d4; 	    wvalid_rom[  165] = 0; 
    i_addr_rom[  166] = 'h00000138; 	    d_addr_rom[  166] = 'h000008d4; 	    wdata_rom[  166] = 'h11587e27; 	    wvalid_rom[  166] = 0; 
    i_addr_rom[  167] = 'h0000074c; 	    d_addr_rom[  167] = 'h00000bf0; 	    wdata_rom[  167] = 'h399a3f3e; 	    wvalid_rom[  167] = 0; 
    i_addr_rom[  168] = 'h00000290; 	    d_addr_rom[  168] = 'h000009ac; 	    wdata_rom[  168] = 'h1eac4642; 	    wvalid_rom[  168] = 1; 
    i_addr_rom[  169] = 'h000005b8; 	    d_addr_rom[  169] = 'h00000c5c; 	    wdata_rom[  169] = 'h079cbb24; 	    wvalid_rom[  169] = 1; 
    i_addr_rom[  170] = 'h00000268; 	    d_addr_rom[  170] = 'h00000e64; 	    wdata_rom[  170] = 'h19faeac7; 	    wvalid_rom[  170] = 0; 
    i_addr_rom[  171] = 'h0000072c; 	    d_addr_rom[  171] = 'h00000dcc; 	    wdata_rom[  171] = 'h716eb1e7; 	    wvalid_rom[  171] = 0; 
    i_addr_rom[  172] = 'h00000540; 	    d_addr_rom[  172] = 'h000009d0; 	    wdata_rom[  172] = 'h3b391c6f; 	    wvalid_rom[  172] = 0; 
    i_addr_rom[  173] = 'h000005c4; 	    d_addr_rom[  173] = 'h00000aa8; 	    wdata_rom[  173] = 'ha0122a28; 	    wvalid_rom[  173] = 1; 
    i_addr_rom[  174] = 'h0000014c; 	    d_addr_rom[  174] = 'h00000bb8; 	    wdata_rom[  174] = 'hda338e3e; 	    wvalid_rom[  174] = 1; 
    i_addr_rom[  175] = 'h00000654; 	    d_addr_rom[  175] = 'h00000950; 	    wdata_rom[  175] = 'h33788ee0; 	    wvalid_rom[  175] = 0; 
    i_addr_rom[  176] = 'h000005a8; 	    d_addr_rom[  176] = 'h00000fbc; 	    wdata_rom[  176] = 'h79b28ad1; 	    wvalid_rom[  176] = 1; 
    i_addr_rom[  177] = 'h000003fc; 	    d_addr_rom[  177] = 'h00000e68; 	    wdata_rom[  177] = 'h20a8b537; 	    wvalid_rom[  177] = 0; 
    i_addr_rom[  178] = 'h00000748; 	    d_addr_rom[  178] = 'h000008a0; 	    wdata_rom[  178] = 'hb9d3828b; 	    wvalid_rom[  178] = 0; 
    i_addr_rom[  179] = 'h000004e8; 	    d_addr_rom[  179] = 'h0000082c; 	    wdata_rom[  179] = 'h92c7bf28; 	    wvalid_rom[  179] = 0; 
    i_addr_rom[  180] = 'h0000022c; 	    d_addr_rom[  180] = 'h00000a1c; 	    wdata_rom[  180] = 'h8db9c6a9; 	    wvalid_rom[  180] = 0; 
    i_addr_rom[  181] = 'h00000454; 	    d_addr_rom[  181] = 'h00000f14; 	    wdata_rom[  181] = 'hfebfc38e; 	    wvalid_rom[  181] = 1; 
    i_addr_rom[  182] = 'h00000064; 	    d_addr_rom[  182] = 'h00000c54; 	    wdata_rom[  182] = 'hd055979f; 	    wvalid_rom[  182] = 1; 
    i_addr_rom[  183] = 'h00000560; 	    d_addr_rom[  183] = 'h000009e8; 	    wdata_rom[  183] = 'h3e59fdaa; 	    wvalid_rom[  183] = 0; 
    i_addr_rom[  184] = 'h00000540; 	    d_addr_rom[  184] = 'h00000b88; 	    wdata_rom[  184] = 'h8a48b06d; 	    wvalid_rom[  184] = 1; 
    i_addr_rom[  185] = 'h0000020c; 	    d_addr_rom[  185] = 'h00000ad0; 	    wdata_rom[  185] = 'h0f3e0e44; 	    wvalid_rom[  185] = 1; 
    i_addr_rom[  186] = 'h00000308; 	    d_addr_rom[  186] = 'h00000e28; 	    wdata_rom[  186] = 'h3b6f207c; 	    wvalid_rom[  186] = 1; 
    i_addr_rom[  187] = 'h000001b4; 	    d_addr_rom[  187] = 'h00000940; 	    wdata_rom[  187] = 'h0e7a70ab; 	    wvalid_rom[  187] = 1; 
    i_addr_rom[  188] = 'h00000350; 	    d_addr_rom[  188] = 'h00000ecc; 	    wdata_rom[  188] = 'h3b2c5df3; 	    wvalid_rom[  188] = 0; 
    i_addr_rom[  189] = 'h00000410; 	    d_addr_rom[  189] = 'h00000bc4; 	    wdata_rom[  189] = 'h108a8745; 	    wvalid_rom[  189] = 1; 
    i_addr_rom[  190] = 'h00000398; 	    d_addr_rom[  190] = 'h0000095c; 	    wdata_rom[  190] = 'hd6af2495; 	    wvalid_rom[  190] = 1; 
    i_addr_rom[  191] = 'h00000728; 	    d_addr_rom[  191] = 'h00000830; 	    wdata_rom[  191] = 'h3917a7eb; 	    wvalid_rom[  191] = 0; 
    i_addr_rom[  192] = 'h00000404; 	    d_addr_rom[  192] = 'h00000b5c; 	    wdata_rom[  192] = 'h74db94a0; 	    wvalid_rom[  192] = 1; 
    i_addr_rom[  193] = 'h00000620; 	    d_addr_rom[  193] = 'h00000e34; 	    wdata_rom[  193] = 'he4e20996; 	    wvalid_rom[  193] = 0; 
    i_addr_rom[  194] = 'h00000798; 	    d_addr_rom[  194] = 'h00000944; 	    wdata_rom[  194] = 'hbac02fe3; 	    wvalid_rom[  194] = 1; 
    i_addr_rom[  195] = 'h000001a0; 	    d_addr_rom[  195] = 'h00000adc; 	    wdata_rom[  195] = 'hae34aff8; 	    wvalid_rom[  195] = 0; 
    i_addr_rom[  196] = 'h00000760; 	    d_addr_rom[  196] = 'h00000b10; 	    wdata_rom[  196] = 'h26bbdd7f; 	    wvalid_rom[  196] = 0; 
    i_addr_rom[  197] = 'h00000624; 	    d_addr_rom[  197] = 'h0000091c; 	    wdata_rom[  197] = 'h538bbd9b; 	    wvalid_rom[  197] = 0; 
    i_addr_rom[  198] = 'h00000368; 	    d_addr_rom[  198] = 'h00000f54; 	    wdata_rom[  198] = 'hce7b4470; 	    wvalid_rom[  198] = 1; 
    i_addr_rom[  199] = 'h00000178; 	    d_addr_rom[  199] = 'h00000e14; 	    wdata_rom[  199] = 'h57e8ae1d; 	    wvalid_rom[  199] = 1; 
    i_addr_rom[  200] = 'h00000000; 	    d_addr_rom[  200] = 'h00000af8; 	    wdata_rom[  200] = 'hcbc3b584; 	    wvalid_rom[  200] = 1; 
    i_addr_rom[  201] = 'h000007f0; 	    d_addr_rom[  201] = 'h00000dc0; 	    wdata_rom[  201] = 'h394ad2e7; 	    wvalid_rom[  201] = 1; 
    i_addr_rom[  202] = 'h000007a8; 	    d_addr_rom[  202] = 'h00000f50; 	    wdata_rom[  202] = 'hc049715f; 	    wvalid_rom[  202] = 1; 
    i_addr_rom[  203] = 'h000000ac; 	    d_addr_rom[  203] = 'h000008ec; 	    wdata_rom[  203] = 'h5738dd27; 	    wvalid_rom[  203] = 1; 
    i_addr_rom[  204] = 'h00000610; 	    d_addr_rom[  204] = 'h00000c34; 	    wdata_rom[  204] = 'h17dec8bd; 	    wvalid_rom[  204] = 0; 
    i_addr_rom[  205] = 'h0000032c; 	    d_addr_rom[  205] = 'h00000a84; 	    wdata_rom[  205] = 'hc1ac49c9; 	    wvalid_rom[  205] = 1; 
    i_addr_rom[  206] = 'h00000674; 	    d_addr_rom[  206] = 'h00000804; 	    wdata_rom[  206] = 'he8417c25; 	    wvalid_rom[  206] = 0; 
    i_addr_rom[  207] = 'h00000568; 	    d_addr_rom[  207] = 'h00000d4c; 	    wdata_rom[  207] = 'h8b930146; 	    wvalid_rom[  207] = 1; 
    i_addr_rom[  208] = 'h00000350; 	    d_addr_rom[  208] = 'h00000db4; 	    wdata_rom[  208] = 'h8149ee66; 	    wvalid_rom[  208] = 1; 
    i_addr_rom[  209] = 'h00000520; 	    d_addr_rom[  209] = 'h00000f88; 	    wdata_rom[  209] = 'hcbeb7477; 	    wvalid_rom[  209] = 0; 
    i_addr_rom[  210] = 'h00000118; 	    d_addr_rom[  210] = 'h00000c9c; 	    wdata_rom[  210] = 'h3444fc97; 	    wvalid_rom[  210] = 0; 
    i_addr_rom[  211] = 'h0000038c; 	    d_addr_rom[  211] = 'h00000ddc; 	    wdata_rom[  211] = 'h33780693; 	    wvalid_rom[  211] = 0; 
    i_addr_rom[  212] = 'h0000053c; 	    d_addr_rom[  212] = 'h0000086c; 	    wdata_rom[  212] = 'h73e3f57e; 	    wvalid_rom[  212] = 1; 
    i_addr_rom[  213] = 'h000002a0; 	    d_addr_rom[  213] = 'h00000c6c; 	    wdata_rom[  213] = 'hd3a60ce9; 	    wvalid_rom[  213] = 0; 
    i_addr_rom[  214] = 'h00000044; 	    d_addr_rom[  214] = 'h00000aac; 	    wdata_rom[  214] = 'h6aaf86ff; 	    wvalid_rom[  214] = 0; 
    i_addr_rom[  215] = 'h00000590; 	    d_addr_rom[  215] = 'h00000e64; 	    wdata_rom[  215] = 'h986627d8; 	    wvalid_rom[  215] = 1; 
    i_addr_rom[  216] = 'h00000590; 	    d_addr_rom[  216] = 'h00000c78; 	    wdata_rom[  216] = 'h9bf7867a; 	    wvalid_rom[  216] = 0; 
    i_addr_rom[  217] = 'h000003ac; 	    d_addr_rom[  217] = 'h00000ef8; 	    wdata_rom[  217] = 'h99a65f93; 	    wvalid_rom[  217] = 1; 
    i_addr_rom[  218] = 'h0000032c; 	    d_addr_rom[  218] = 'h00000e4c; 	    wdata_rom[  218] = 'h04d95a34; 	    wvalid_rom[  218] = 0; 
    i_addr_rom[  219] = 'h00000168; 	    d_addr_rom[  219] = 'h0000094c; 	    wdata_rom[  219] = 'hd0bebcbe; 	    wvalid_rom[  219] = 0; 
    i_addr_rom[  220] = 'h00000444; 	    d_addr_rom[  220] = 'h00000bf8; 	    wdata_rom[  220] = 'hf977a14b; 	    wvalid_rom[  220] = 1; 
    i_addr_rom[  221] = 'h0000021c; 	    d_addr_rom[  221] = 'h00000ce0; 	    wdata_rom[  221] = 'h39cbeb94; 	    wvalid_rom[  221] = 1; 
    i_addr_rom[  222] = 'h000005b0; 	    d_addr_rom[  222] = 'h00000c1c; 	    wdata_rom[  222] = 'h0d64f941; 	    wvalid_rom[  222] = 0; 
    i_addr_rom[  223] = 'h000000a8; 	    d_addr_rom[  223] = 'h000008e4; 	    wdata_rom[  223] = 'h9ccdd8e2; 	    wvalid_rom[  223] = 1; 
    i_addr_rom[  224] = 'h0000052c; 	    d_addr_rom[  224] = 'h00000b7c; 	    wdata_rom[  224] = 'hb87b66be; 	    wvalid_rom[  224] = 1; 
    i_addr_rom[  225] = 'h000007ac; 	    d_addr_rom[  225] = 'h00000c60; 	    wdata_rom[  225] = 'h98881585; 	    wvalid_rom[  225] = 1; 
    i_addr_rom[  226] = 'h000003fc; 	    d_addr_rom[  226] = 'h00000840; 	    wdata_rom[  226] = 'h71dd29e7; 	    wvalid_rom[  226] = 1; 
    i_addr_rom[  227] = 'h00000574; 	    d_addr_rom[  227] = 'h00000b4c; 	    wdata_rom[  227] = 'h5b69538b; 	    wvalid_rom[  227] = 1; 
    i_addr_rom[  228] = 'h00000530; 	    d_addr_rom[  228] = 'h00000e14; 	    wdata_rom[  228] = 'h2fd69a70; 	    wvalid_rom[  228] = 0; 
    i_addr_rom[  229] = 'h00000628; 	    d_addr_rom[  229] = 'h00000f84; 	    wdata_rom[  229] = 'h1bde1ea0; 	    wvalid_rom[  229] = 0; 
    i_addr_rom[  230] = 'h00000340; 	    d_addr_rom[  230] = 'h000008f4; 	    wdata_rom[  230] = 'h86c234e4; 	    wvalid_rom[  230] = 1; 
    i_addr_rom[  231] = 'h000003e0; 	    d_addr_rom[  231] = 'h00000c00; 	    wdata_rom[  231] = 'h1833b2d6; 	    wvalid_rom[  231] = 0; 
    i_addr_rom[  232] = 'h00000574; 	    d_addr_rom[  232] = 'h00000cd8; 	    wdata_rom[  232] = 'hb007d04d; 	    wvalid_rom[  232] = 1; 
    i_addr_rom[  233] = 'h0000061c; 	    d_addr_rom[  233] = 'h00000b14; 	    wdata_rom[  233] = 'h9747c5e9; 	    wvalid_rom[  233] = 1; 
    i_addr_rom[  234] = 'h00000328; 	    d_addr_rom[  234] = 'h00000ca4; 	    wdata_rom[  234] = 'h4c5d3cc9; 	    wvalid_rom[  234] = 0; 
    i_addr_rom[  235] = 'h00000140; 	    d_addr_rom[  235] = 'h00000e18; 	    wdata_rom[  235] = 'hfecd6d5b; 	    wvalid_rom[  235] = 0; 
    i_addr_rom[  236] = 'h00000668; 	    d_addr_rom[  236] = 'h00000c7c; 	    wdata_rom[  236] = 'h6a975fc5; 	    wvalid_rom[  236] = 0; 
    i_addr_rom[  237] = 'h000001c4; 	    d_addr_rom[  237] = 'h000008e8; 	    wdata_rom[  237] = 'hfe87adbf; 	    wvalid_rom[  237] = 0; 
    i_addr_rom[  238] = 'h000006dc; 	    d_addr_rom[  238] = 'h00000abc; 	    wdata_rom[  238] = 'hd2586ea2; 	    wvalid_rom[  238] = 1; 
    i_addr_rom[  239] = 'h000000b4; 	    d_addr_rom[  239] = 'h00000a88; 	    wdata_rom[  239] = 'h3be1791b; 	    wvalid_rom[  239] = 0; 
    i_addr_rom[  240] = 'h000004bc; 	    d_addr_rom[  240] = 'h0000092c; 	    wdata_rom[  240] = 'h7c589062; 	    wvalid_rom[  240] = 1; 
    i_addr_rom[  241] = 'h00000708; 	    d_addr_rom[  241] = 'h00000bb0; 	    wdata_rom[  241] = 'ha25825fb; 	    wvalid_rom[  241] = 1; 
    i_addr_rom[  242] = 'h000005dc; 	    d_addr_rom[  242] = 'h00000fa4; 	    wdata_rom[  242] = 'he2f599c5; 	    wvalid_rom[  242] = 0; 
    i_addr_rom[  243] = 'h00000280; 	    d_addr_rom[  243] = 'h00000a9c; 	    wdata_rom[  243] = 'hcea6089e; 	    wvalid_rom[  243] = 0; 
    i_addr_rom[  244] = 'h0000072c; 	    d_addr_rom[  244] = 'h00000c4c; 	    wdata_rom[  244] = 'hbfc91d77; 	    wvalid_rom[  244] = 1; 
    i_addr_rom[  245] = 'h000002fc; 	    d_addr_rom[  245] = 'h00000dd4; 	    wdata_rom[  245] = 'h4429d10b; 	    wvalid_rom[  245] = 0; 
    i_addr_rom[  246] = 'h000005f4; 	    d_addr_rom[  246] = 'h00000fb4; 	    wdata_rom[  246] = 'h7e68b1a3; 	    wvalid_rom[  246] = 1; 
    i_addr_rom[  247] = 'h0000077c; 	    d_addr_rom[  247] = 'h000008d0; 	    wdata_rom[  247] = 'h491b130e; 	    wvalid_rom[  247] = 0; 
    i_addr_rom[  248] = 'h00000228; 	    d_addr_rom[  248] = 'h00000af4; 	    wdata_rom[  248] = 'hebd356b9; 	    wvalid_rom[  248] = 0; 
    i_addr_rom[  249] = 'h00000664; 	    d_addr_rom[  249] = 'h00000d40; 	    wdata_rom[  249] = 'haa0b1ff7; 	    wvalid_rom[  249] = 1; 
    i_addr_rom[  250] = 'h00000748; 	    d_addr_rom[  250] = 'h00000ee8; 	    wdata_rom[  250] = 'h1cdf8595; 	    wvalid_rom[  250] = 0; 
    i_addr_rom[  251] = 'h00000198; 	    d_addr_rom[  251] = 'h00000b90; 	    wdata_rom[  251] = 'h63bbb0ba; 	    wvalid_rom[  251] = 0; 
    i_addr_rom[  252] = 'h00000254; 	    d_addr_rom[  252] = 'h00000f90; 	    wdata_rom[  252] = 'h48305f63; 	    wvalid_rom[  252] = 0; 
    i_addr_rom[  253] = 'h00000100; 	    d_addr_rom[  253] = 'h00000fb8; 	    wdata_rom[  253] = 'h1f790323; 	    wvalid_rom[  253] = 1; 
    i_addr_rom[  254] = 'h000007b4; 	    d_addr_rom[  254] = 'h00000c04; 	    wdata_rom[  254] = 'haef4ad49; 	    wvalid_rom[  254] = 0; 
    i_addr_rom[  255] = 'h00000780; 	    d_addr_rom[  255] = 'h00000db0; 	    wdata_rom[  255] = 'h74167e10; 	    wvalid_rom[  255] = 0; 
    i_addr_rom[  256] = 'h0000072c; 	    d_addr_rom[  256] = 'h00000e6c; 	    wdata_rom[  256] = 'h1dd690c8; 	    wvalid_rom[  256] = 0; 
    i_addr_rom[  257] = 'h00000520; 	    d_addr_rom[  257] = 'h0000096c; 	    wdata_rom[  257] = 'h13b2d19a; 	    wvalid_rom[  257] = 1; 
    i_addr_rom[  258] = 'h00000714; 	    d_addr_rom[  258] = 'h00000c20; 	    wdata_rom[  258] = 'hd07a13da; 	    wvalid_rom[  258] = 0; 
    i_addr_rom[  259] = 'h00000248; 	    d_addr_rom[  259] = 'h00000acc; 	    wdata_rom[  259] = 'hf1627121; 	    wvalid_rom[  259] = 1; 
    i_addr_rom[  260] = 'h000005e4; 	    d_addr_rom[  260] = 'h00000c3c; 	    wdata_rom[  260] = 'h4ff30713; 	    wvalid_rom[  260] = 0; 
    i_addr_rom[  261] = 'h000006d8; 	    d_addr_rom[  261] = 'h00000b1c; 	    wdata_rom[  261] = 'hc22ffe69; 	    wvalid_rom[  261] = 1; 
    i_addr_rom[  262] = 'h00000188; 	    d_addr_rom[  262] = 'h00000e7c; 	    wdata_rom[  262] = 'he4b7bb92; 	    wvalid_rom[  262] = 0; 
    i_addr_rom[  263] = 'h00000410; 	    d_addr_rom[  263] = 'h00000930; 	    wdata_rom[  263] = 'h35bb7191; 	    wvalid_rom[  263] = 1; 
    i_addr_rom[  264] = 'h000004e0; 	    d_addr_rom[  264] = 'h00000ed4; 	    wdata_rom[  264] = 'hf7bdd3a2; 	    wvalid_rom[  264] = 0; 
    i_addr_rom[  265] = 'h000004a8; 	    d_addr_rom[  265] = 'h00000ad4; 	    wdata_rom[  265] = 'hd7bc4679; 	    wvalid_rom[  265] = 0; 
    i_addr_rom[  266] = 'h00000628; 	    d_addr_rom[  266] = 'h00000c3c; 	    wdata_rom[  266] = 'ha1b2dfa9; 	    wvalid_rom[  266] = 1; 
    i_addr_rom[  267] = 'h00000480; 	    d_addr_rom[  267] = 'h00000f10; 	    wdata_rom[  267] = 'h3dc0704b; 	    wvalid_rom[  267] = 0; 
    i_addr_rom[  268] = 'h00000538; 	    d_addr_rom[  268] = 'h00000afc; 	    wdata_rom[  268] = 'hb3ca3ea9; 	    wvalid_rom[  268] = 1; 
    i_addr_rom[  269] = 'h00000270; 	    d_addr_rom[  269] = 'h00000a54; 	    wdata_rom[  269] = 'hd6d142c6; 	    wvalid_rom[  269] = 1; 
    i_addr_rom[  270] = 'h00000104; 	    d_addr_rom[  270] = 'h0000087c; 	    wdata_rom[  270] = 'hc7375594; 	    wvalid_rom[  270] = 0; 
    i_addr_rom[  271] = 'h00000350; 	    d_addr_rom[  271] = 'h00000d04; 	    wdata_rom[  271] = 'h7dcff8d9; 	    wvalid_rom[  271] = 0; 
    i_addr_rom[  272] = 'h00000684; 	    d_addr_rom[  272] = 'h00000fc8; 	    wdata_rom[  272] = 'h85e02a93; 	    wvalid_rom[  272] = 0; 
    i_addr_rom[  273] = 'h00000210; 	    d_addr_rom[  273] = 'h00000f3c; 	    wdata_rom[  273] = 'hdd8c6062; 	    wvalid_rom[  273] = 0; 
    i_addr_rom[  274] = 'h0000043c; 	    d_addr_rom[  274] = 'h00000fec; 	    wdata_rom[  274] = 'h5f64b6a2; 	    wvalid_rom[  274] = 1; 
    i_addr_rom[  275] = 'h00000720; 	    d_addr_rom[  275] = 'h00000ff8; 	    wdata_rom[  275] = 'hf3eec535; 	    wvalid_rom[  275] = 0; 
    i_addr_rom[  276] = 'h00000180; 	    d_addr_rom[  276] = 'h00000bd4; 	    wdata_rom[  276] = 'h3b2c4614; 	    wvalid_rom[  276] = 1; 
    i_addr_rom[  277] = 'h000003e8; 	    d_addr_rom[  277] = 'h00000fc8; 	    wdata_rom[  277] = 'h834f5279; 	    wvalid_rom[  277] = 1; 
    i_addr_rom[  278] = 'h000003a8; 	    d_addr_rom[  278] = 'h00000fc8; 	    wdata_rom[  278] = 'h2d6b83d9; 	    wvalid_rom[  278] = 1; 
    i_addr_rom[  279] = 'h000005e4; 	    d_addr_rom[  279] = 'h00000974; 	    wdata_rom[  279] = 'he42eedb3; 	    wvalid_rom[  279] = 1; 
    i_addr_rom[  280] = 'h00000280; 	    d_addr_rom[  280] = 'h00000b28; 	    wdata_rom[  280] = 'hf4030983; 	    wvalid_rom[  280] = 0; 
    i_addr_rom[  281] = 'h000006b4; 	    d_addr_rom[  281] = 'h00000c0c; 	    wdata_rom[  281] = 'hcb4e211c; 	    wvalid_rom[  281] = 1; 
    i_addr_rom[  282] = 'h000005c8; 	    d_addr_rom[  282] = 'h00000e90; 	    wdata_rom[  282] = 'hf5d2b767; 	    wvalid_rom[  282] = 0; 
    i_addr_rom[  283] = 'h00000208; 	    d_addr_rom[  283] = 'h000008cc; 	    wdata_rom[  283] = 'h60e3efd2; 	    wvalid_rom[  283] = 1; 
    i_addr_rom[  284] = 'h00000228; 	    d_addr_rom[  284] = 'h00000bb0; 	    wdata_rom[  284] = 'hf7bfef83; 	    wvalid_rom[  284] = 0; 
    i_addr_rom[  285] = 'h000004e0; 	    d_addr_rom[  285] = 'h00000c70; 	    wdata_rom[  285] = 'h66ac85cd; 	    wvalid_rom[  285] = 0; 
    i_addr_rom[  286] = 'h000003ec; 	    d_addr_rom[  286] = 'h00000900; 	    wdata_rom[  286] = 'h14f72a39; 	    wvalid_rom[  286] = 1; 
    i_addr_rom[  287] = 'h00000628; 	    d_addr_rom[  287] = 'h00000ee0; 	    wdata_rom[  287] = 'h7d85d31f; 	    wvalid_rom[  287] = 0; 
    i_addr_rom[  288] = 'h000002e4; 	    d_addr_rom[  288] = 'h00000dd8; 	    wdata_rom[  288] = 'haac02c86; 	    wvalid_rom[  288] = 1; 
    i_addr_rom[  289] = 'h000000ac; 	    d_addr_rom[  289] = 'h00000f9c; 	    wdata_rom[  289] = 'ha8cde139; 	    wvalid_rom[  289] = 1; 
    i_addr_rom[  290] = 'h00000170; 	    d_addr_rom[  290] = 'h00000ee4; 	    wdata_rom[  290] = 'h41989dbf; 	    wvalid_rom[  290] = 0; 
    i_addr_rom[  291] = 'h00000794; 	    d_addr_rom[  291] = 'h00000a20; 	    wdata_rom[  291] = 'h87e574bb; 	    wvalid_rom[  291] = 1; 
    i_addr_rom[  292] = 'h000005ac; 	    d_addr_rom[  292] = 'h00000f68; 	    wdata_rom[  292] = 'h8b750863; 	    wvalid_rom[  292] = 1; 
    i_addr_rom[  293] = 'h0000036c; 	    d_addr_rom[  293] = 'h00000de0; 	    wdata_rom[  293] = 'hc64e1925; 	    wvalid_rom[  293] = 1; 
    i_addr_rom[  294] = 'h0000072c; 	    d_addr_rom[  294] = 'h000009f0; 	    wdata_rom[  294] = 'hedd351a3; 	    wvalid_rom[  294] = 1; 
    i_addr_rom[  295] = 'h0000007c; 	    d_addr_rom[  295] = 'h00000adc; 	    wdata_rom[  295] = 'h4f70d02b; 	    wvalid_rom[  295] = 1; 
    i_addr_rom[  296] = 'h00000188; 	    d_addr_rom[  296] = 'h00000cc4; 	    wdata_rom[  296] = 'hb9892927; 	    wvalid_rom[  296] = 0; 
    i_addr_rom[  297] = 'h00000758; 	    d_addr_rom[  297] = 'h00000f98; 	    wdata_rom[  297] = 'hb0817a5b; 	    wvalid_rom[  297] = 1; 
    i_addr_rom[  298] = 'h00000100; 	    d_addr_rom[  298] = 'h00000d7c; 	    wdata_rom[  298] = 'hb34a45a5; 	    wvalid_rom[  298] = 0; 
    i_addr_rom[  299] = 'h000006b8; 	    d_addr_rom[  299] = 'h00000b20; 	    wdata_rom[  299] = 'h19047fe3; 	    wvalid_rom[  299] = 0; 
    i_addr_rom[  300] = 'h0000015c; 	    d_addr_rom[  300] = 'h00000ed0; 	    wdata_rom[  300] = 'haeb5e66c; 	    wvalid_rom[  300] = 0; 
    i_addr_rom[  301] = 'h00000608; 	    d_addr_rom[  301] = 'h00000954; 	    wdata_rom[  301] = 'hc2c313ef; 	    wvalid_rom[  301] = 1; 
    i_addr_rom[  302] = 'h000007c0; 	    d_addr_rom[  302] = 'h00000d60; 	    wdata_rom[  302] = 'hc22bf88f; 	    wvalid_rom[  302] = 0; 
    i_addr_rom[  303] = 'h0000023c; 	    d_addr_rom[  303] = 'h00000aac; 	    wdata_rom[  303] = 'h1ba73471; 	    wvalid_rom[  303] = 0; 
    i_addr_rom[  304] = 'h00000250; 	    d_addr_rom[  304] = 'h00000dac; 	    wdata_rom[  304] = 'h1d2b9594; 	    wvalid_rom[  304] = 0; 
    i_addr_rom[  305] = 'h000003e4; 	    d_addr_rom[  305] = 'h00000a70; 	    wdata_rom[  305] = 'h8c6a52f2; 	    wvalid_rom[  305] = 1; 
    i_addr_rom[  306] = 'h00000778; 	    d_addr_rom[  306] = 'h00000820; 	    wdata_rom[  306] = 'h39ba9990; 	    wvalid_rom[  306] = 0; 
    i_addr_rom[  307] = 'h000004f8; 	    d_addr_rom[  307] = 'h00000fcc; 	    wdata_rom[  307] = 'h8c12bd26; 	    wvalid_rom[  307] = 1; 
    i_addr_rom[  308] = 'h0000010c; 	    d_addr_rom[  308] = 'h00000cb4; 	    wdata_rom[  308] = 'h915b252c; 	    wvalid_rom[  308] = 1; 
    i_addr_rom[  309] = 'h0000066c; 	    d_addr_rom[  309] = 'h00000cc0; 	    wdata_rom[  309] = 'h44a75845; 	    wvalid_rom[  309] = 1; 
    i_addr_rom[  310] = 'h000005cc; 	    d_addr_rom[  310] = 'h00000b5c; 	    wdata_rom[  310] = 'ha1d66459; 	    wvalid_rom[  310] = 0; 
    i_addr_rom[  311] = 'h000000a4; 	    d_addr_rom[  311] = 'h00000bbc; 	    wdata_rom[  311] = 'hff132cd4; 	    wvalid_rom[  311] = 0; 
    i_addr_rom[  312] = 'h00000374; 	    d_addr_rom[  312] = 'h00000b70; 	    wdata_rom[  312] = 'h737ea78d; 	    wvalid_rom[  312] = 0; 
    i_addr_rom[  313] = 'h000006f8; 	    d_addr_rom[  313] = 'h00000e04; 	    wdata_rom[  313] = 'h46614d16; 	    wvalid_rom[  313] = 0; 
    i_addr_rom[  314] = 'h000006c4; 	    d_addr_rom[  314] = 'h00000b8c; 	    wdata_rom[  314] = 'h2253c33f; 	    wvalid_rom[  314] = 1; 
    i_addr_rom[  315] = 'h00000148; 	    d_addr_rom[  315] = 'h00000a38; 	    wdata_rom[  315] = 'hbf393f30; 	    wvalid_rom[  315] = 1; 
    i_addr_rom[  316] = 'h00000388; 	    d_addr_rom[  316] = 'h00000c3c; 	    wdata_rom[  316] = 'hea511a3a; 	    wvalid_rom[  316] = 1; 
    i_addr_rom[  317] = 'h0000020c; 	    d_addr_rom[  317] = 'h00000a84; 	    wdata_rom[  317] = 'h6916578f; 	    wvalid_rom[  317] = 1; 
    i_addr_rom[  318] = 'h00000388; 	    d_addr_rom[  318] = 'h00000d7c; 	    wdata_rom[  318] = 'h3aa1690a; 	    wvalid_rom[  318] = 1; 
    i_addr_rom[  319] = 'h00000308; 	    d_addr_rom[  319] = 'h00000b18; 	    wdata_rom[  319] = 'hb40db2fa; 	    wvalid_rom[  319] = 0; 
    i_addr_rom[  320] = 'h000001f0; 	    d_addr_rom[  320] = 'h00000ebc; 	    wdata_rom[  320] = 'h56ce7bf6; 	    wvalid_rom[  320] = 0; 
    i_addr_rom[  321] = 'h000007a4; 	    d_addr_rom[  321] = 'h00000a70; 	    wdata_rom[  321] = 'h5b0a1bb7; 	    wvalid_rom[  321] = 0; 
    i_addr_rom[  322] = 'h00000280; 	    d_addr_rom[  322] = 'h00000c60; 	    wdata_rom[  322] = 'h3d6c3358; 	    wvalid_rom[  322] = 0; 
    i_addr_rom[  323] = 'h0000026c; 	    d_addr_rom[  323] = 'h00000f94; 	    wdata_rom[  323] = 'h0a1ae027; 	    wvalid_rom[  323] = 1; 
    i_addr_rom[  324] = 'h000004b4; 	    d_addr_rom[  324] = 'h00000c18; 	    wdata_rom[  324] = 'h4c62aaab; 	    wvalid_rom[  324] = 0; 
    i_addr_rom[  325] = 'h000005b4; 	    d_addr_rom[  325] = 'h000008a0; 	    wdata_rom[  325] = 'h64e89eec; 	    wvalid_rom[  325] = 0; 
    i_addr_rom[  326] = 'h00000594; 	    d_addr_rom[  326] = 'h00000e04; 	    wdata_rom[  326] = 'he52b725f; 	    wvalid_rom[  326] = 0; 
    i_addr_rom[  327] = 'h000005dc; 	    d_addr_rom[  327] = 'h00000a78; 	    wdata_rom[  327] = 'he49ee69a; 	    wvalid_rom[  327] = 0; 
    i_addr_rom[  328] = 'h000001ac; 	    d_addr_rom[  328] = 'h00000f84; 	    wdata_rom[  328] = 'hea30e483; 	    wvalid_rom[  328] = 0; 
    i_addr_rom[  329] = 'h000007d4; 	    d_addr_rom[  329] = 'h00000cd4; 	    wdata_rom[  329] = 'hf2880d70; 	    wvalid_rom[  329] = 0; 
    i_addr_rom[  330] = 'h00000740; 	    d_addr_rom[  330] = 'h00000d34; 	    wdata_rom[  330] = 'h3360f233; 	    wvalid_rom[  330] = 1; 
    i_addr_rom[  331] = 'h000007e0; 	    d_addr_rom[  331] = 'h00000fa4; 	    wdata_rom[  331] = 'hfa3451ca; 	    wvalid_rom[  331] = 0; 
    i_addr_rom[  332] = 'h00000598; 	    d_addr_rom[  332] = 'h00000ab8; 	    wdata_rom[  332] = 'hf71602e8; 	    wvalid_rom[  332] = 0; 
    i_addr_rom[  333] = 'h000000d4; 	    d_addr_rom[  333] = 'h00000998; 	    wdata_rom[  333] = 'h96a4342c; 	    wvalid_rom[  333] = 0; 
    i_addr_rom[  334] = 'h000001d0; 	    d_addr_rom[  334] = 'h00000fe8; 	    wdata_rom[  334] = 'h8aadd95f; 	    wvalid_rom[  334] = 0; 
    i_addr_rom[  335] = 'h00000530; 	    d_addr_rom[  335] = 'h00000bfc; 	    wdata_rom[  335] = 'h100e49c7; 	    wvalid_rom[  335] = 1; 
    i_addr_rom[  336] = 'h000002c8; 	    d_addr_rom[  336] = 'h00000bc8; 	    wdata_rom[  336] = 'he853d7f2; 	    wvalid_rom[  336] = 0; 
    i_addr_rom[  337] = 'h000006e0; 	    d_addr_rom[  337] = 'h0000091c; 	    wdata_rom[  337] = 'h27965579; 	    wvalid_rom[  337] = 1; 
    i_addr_rom[  338] = 'h00000038; 	    d_addr_rom[  338] = 'h00000820; 	    wdata_rom[  338] = 'h9192227b; 	    wvalid_rom[  338] = 0; 
    i_addr_rom[  339] = 'h0000062c; 	    d_addr_rom[  339] = 'h00000eb0; 	    wdata_rom[  339] = 'hdc697929; 	    wvalid_rom[  339] = 1; 
    i_addr_rom[  340] = 'h000004e8; 	    d_addr_rom[  340] = 'h00000db4; 	    wdata_rom[  340] = 'h95313a48; 	    wvalid_rom[  340] = 1; 
    i_addr_rom[  341] = 'h00000640; 	    d_addr_rom[  341] = 'h00000c9c; 	    wdata_rom[  341] = 'hd55d418e; 	    wvalid_rom[  341] = 0; 
    i_addr_rom[  342] = 'h000001cc; 	    d_addr_rom[  342] = 'h00000d38; 	    wdata_rom[  342] = 'ha3a73f0d; 	    wvalid_rom[  342] = 0; 
    i_addr_rom[  343] = 'h000005bc; 	    d_addr_rom[  343] = 'h00000bf8; 	    wdata_rom[  343] = 'h964e7502; 	    wvalid_rom[  343] = 0; 
    i_addr_rom[  344] = 'h00000178; 	    d_addr_rom[  344] = 'h00000d68; 	    wdata_rom[  344] = 'h79884e39; 	    wvalid_rom[  344] = 1; 
    i_addr_rom[  345] = 'h00000670; 	    d_addr_rom[  345] = 'h00000da8; 	    wdata_rom[  345] = 'he11b60b7; 	    wvalid_rom[  345] = 1; 
    i_addr_rom[  346] = 'h000000c4; 	    d_addr_rom[  346] = 'h00000934; 	    wdata_rom[  346] = 'hf76b4442; 	    wvalid_rom[  346] = 1; 
    i_addr_rom[  347] = 'h0000016c; 	    d_addr_rom[  347] = 'h00000ad4; 	    wdata_rom[  347] = 'hc7c8c4eb; 	    wvalid_rom[  347] = 0; 
    i_addr_rom[  348] = 'h00000014; 	    d_addr_rom[  348] = 'h00000f68; 	    wdata_rom[  348] = 'h53c414c4; 	    wvalid_rom[  348] = 0; 
    i_addr_rom[  349] = 'h000007cc; 	    d_addr_rom[  349] = 'h00000acc; 	    wdata_rom[  349] = 'he5f4e61b; 	    wvalid_rom[  349] = 0; 
    i_addr_rom[  350] = 'h000001ec; 	    d_addr_rom[  350] = 'h00000b20; 	    wdata_rom[  350] = 'hb7837603; 	    wvalid_rom[  350] = 0; 
    i_addr_rom[  351] = 'h0000043c; 	    d_addr_rom[  351] = 'h00000e94; 	    wdata_rom[  351] = 'h6eb0e5ad; 	    wvalid_rom[  351] = 1; 
    i_addr_rom[  352] = 'h0000047c; 	    d_addr_rom[  352] = 'h000008dc; 	    wdata_rom[  352] = 'hce610854; 	    wvalid_rom[  352] = 0; 
    i_addr_rom[  353] = 'h0000073c; 	    d_addr_rom[  353] = 'h00000c94; 	    wdata_rom[  353] = 'h18f2a068; 	    wvalid_rom[  353] = 1; 
    i_addr_rom[  354] = 'h000004ac; 	    d_addr_rom[  354] = 'h00000af8; 	    wdata_rom[  354] = 'h3cfc56fb; 	    wvalid_rom[  354] = 1; 
    i_addr_rom[  355] = 'h00000034; 	    d_addr_rom[  355] = 'h00000fbc; 	    wdata_rom[  355] = 'h787748cb; 	    wvalid_rom[  355] = 1; 
    i_addr_rom[  356] = 'h00000768; 	    d_addr_rom[  356] = 'h00000e70; 	    wdata_rom[  356] = 'h6ad7a888; 	    wvalid_rom[  356] = 0; 
    i_addr_rom[  357] = 'h00000764; 	    d_addr_rom[  357] = 'h00000fc4; 	    wdata_rom[  357] = 'h9dc437c9; 	    wvalid_rom[  357] = 0; 
    i_addr_rom[  358] = 'h000007d4; 	    d_addr_rom[  358] = 'h00000d2c; 	    wdata_rom[  358] = 'h24182843; 	    wvalid_rom[  358] = 0; 
    i_addr_rom[  359] = 'h000004cc; 	    d_addr_rom[  359] = 'h00000efc; 	    wdata_rom[  359] = 'h7efaad77; 	    wvalid_rom[  359] = 0; 
    i_addr_rom[  360] = 'h000000a8; 	    d_addr_rom[  360] = 'h00000da4; 	    wdata_rom[  360] = 'hcda27a2e; 	    wvalid_rom[  360] = 0; 
    i_addr_rom[  361] = 'h00000650; 	    d_addr_rom[  361] = 'h000008e8; 	    wdata_rom[  361] = 'h6a5747d1; 	    wvalid_rom[  361] = 1; 
    i_addr_rom[  362] = 'h00000614; 	    d_addr_rom[  362] = 'h00000bac; 	    wdata_rom[  362] = 'hcee61da9; 	    wvalid_rom[  362] = 0; 
    i_addr_rom[  363] = 'h000006fc; 	    d_addr_rom[  363] = 'h00000e3c; 	    wdata_rom[  363] = 'h7eb12fb6; 	    wvalid_rom[  363] = 1; 
    i_addr_rom[  364] = 'h000000a4; 	    d_addr_rom[  364] = 'h000009e8; 	    wdata_rom[  364] = 'hd96519ff; 	    wvalid_rom[  364] = 0; 
    i_addr_rom[  365] = 'h0000051c; 	    d_addr_rom[  365] = 'h000009fc; 	    wdata_rom[  365] = 'h95cf30f5; 	    wvalid_rom[  365] = 1; 
    i_addr_rom[  366] = 'h00000594; 	    d_addr_rom[  366] = 'h00000bdc; 	    wdata_rom[  366] = 'hd421a9dd; 	    wvalid_rom[  366] = 1; 
    i_addr_rom[  367] = 'h000005cc; 	    d_addr_rom[  367] = 'h000008e4; 	    wdata_rom[  367] = 'h4407949e; 	    wvalid_rom[  367] = 1; 
    i_addr_rom[  368] = 'h000003d0; 	    d_addr_rom[  368] = 'h00000860; 	    wdata_rom[  368] = 'h5f0bbc37; 	    wvalid_rom[  368] = 1; 
    i_addr_rom[  369] = 'h00000200; 	    d_addr_rom[  369] = 'h00000a38; 	    wdata_rom[  369] = 'hd08fa385; 	    wvalid_rom[  369] = 1; 
    i_addr_rom[  370] = 'h000001a4; 	    d_addr_rom[  370] = 'h00000d10; 	    wdata_rom[  370] = 'h52100783; 	    wvalid_rom[  370] = 0; 
    i_addr_rom[  371] = 'h00000368; 	    d_addr_rom[  371] = 'h00000980; 	    wdata_rom[  371] = 'hc59ad40f; 	    wvalid_rom[  371] = 0; 
    i_addr_rom[  372] = 'h00000004; 	    d_addr_rom[  372] = 'h00000fb0; 	    wdata_rom[  372] = 'h771eb684; 	    wvalid_rom[  372] = 0; 
    i_addr_rom[  373] = 'h00000588; 	    d_addr_rom[  373] = 'h00000da8; 	    wdata_rom[  373] = 'h114eec15; 	    wvalid_rom[  373] = 1; 
    i_addr_rom[  374] = 'h00000620; 	    d_addr_rom[  374] = 'h00000904; 	    wdata_rom[  374] = 'h15956394; 	    wvalid_rom[  374] = 0; 
    i_addr_rom[  375] = 'h000000c0; 	    d_addr_rom[  375] = 'h00000934; 	    wdata_rom[  375] = 'h9e3bdad5; 	    wvalid_rom[  375] = 1; 
    i_addr_rom[  376] = 'h000002c4; 	    d_addr_rom[  376] = 'h00000fb8; 	    wdata_rom[  376] = 'hb48b890f; 	    wvalid_rom[  376] = 1; 
    i_addr_rom[  377] = 'h000007f4; 	    d_addr_rom[  377] = 'h0000085c; 	    wdata_rom[  377] = 'h34069fde; 	    wvalid_rom[  377] = 0; 
    i_addr_rom[  378] = 'h000000dc; 	    d_addr_rom[  378] = 'h000009c4; 	    wdata_rom[  378] = 'h616a59d7; 	    wvalid_rom[  378] = 1; 
    i_addr_rom[  379] = 'h0000008c; 	    d_addr_rom[  379] = 'h00000fcc; 	    wdata_rom[  379] = 'he17373ad; 	    wvalid_rom[  379] = 1; 
    i_addr_rom[  380] = 'h000006a8; 	    d_addr_rom[  380] = 'h00000bf0; 	    wdata_rom[  380] = 'h203fb171; 	    wvalid_rom[  380] = 1; 
    i_addr_rom[  381] = 'h000002e0; 	    d_addr_rom[  381] = 'h00000cbc; 	    wdata_rom[  381] = 'he8a7fb31; 	    wvalid_rom[  381] = 0; 
    i_addr_rom[  382] = 'h000003e0; 	    d_addr_rom[  382] = 'h00000f38; 	    wdata_rom[  382] = 'h01592ecd; 	    wvalid_rom[  382] = 1; 
    i_addr_rom[  383] = 'h00000760; 	    d_addr_rom[  383] = 'h00000a74; 	    wdata_rom[  383] = 'h04d719d6; 	    wvalid_rom[  383] = 0; 
    i_addr_rom[  384] = 'h0000053c; 	    d_addr_rom[  384] = 'h00000970; 	    wdata_rom[  384] = 'hd56ce797; 	    wvalid_rom[  384] = 0; 
    i_addr_rom[  385] = 'h00000644; 	    d_addr_rom[  385] = 'h00000980; 	    wdata_rom[  385] = 'h928bb4d7; 	    wvalid_rom[  385] = 1; 
    i_addr_rom[  386] = 'h000000f4; 	    d_addr_rom[  386] = 'h00000970; 	    wdata_rom[  386] = 'hcc6bfc42; 	    wvalid_rom[  386] = 1; 
    i_addr_rom[  387] = 'h000007bc; 	    d_addr_rom[  387] = 'h00000f2c; 	    wdata_rom[  387] = 'h9465cfed; 	    wvalid_rom[  387] = 1; 
    i_addr_rom[  388] = 'h00000198; 	    d_addr_rom[  388] = 'h00000f98; 	    wdata_rom[  388] = 'h2ae42015; 	    wvalid_rom[  388] = 0; 
    i_addr_rom[  389] = 'h0000048c; 	    d_addr_rom[  389] = 'h00000984; 	    wdata_rom[  389] = 'hac85d5ca; 	    wvalid_rom[  389] = 1; 
    i_addr_rom[  390] = 'h00000238; 	    d_addr_rom[  390] = 'h00000bcc; 	    wdata_rom[  390] = 'h8b928712; 	    wvalid_rom[  390] = 0; 
    i_addr_rom[  391] = 'h000001d0; 	    d_addr_rom[  391] = 'h00000e38; 	    wdata_rom[  391] = 'h5bc2f6f1; 	    wvalid_rom[  391] = 1; 
    i_addr_rom[  392] = 'h0000021c; 	    d_addr_rom[  392] = 'h00000f68; 	    wdata_rom[  392] = 'h773ca05d; 	    wvalid_rom[  392] = 1; 
    i_addr_rom[  393] = 'h00000720; 	    d_addr_rom[  393] = 'h000008ec; 	    wdata_rom[  393] = 'h94a4af86; 	    wvalid_rom[  393] = 1; 
    i_addr_rom[  394] = 'h00000390; 	    d_addr_rom[  394] = 'h000008ec; 	    wdata_rom[  394] = 'hfad84b80; 	    wvalid_rom[  394] = 0; 
    i_addr_rom[  395] = 'h000005b4; 	    d_addr_rom[  395] = 'h00000dac; 	    wdata_rom[  395] = 'hf7e2f71a; 	    wvalid_rom[  395] = 1; 
    i_addr_rom[  396] = 'h00000310; 	    d_addr_rom[  396] = 'h00000cd8; 	    wdata_rom[  396] = 'hb80a08ea; 	    wvalid_rom[  396] = 1; 
    i_addr_rom[  397] = 'h000000b4; 	    d_addr_rom[  397] = 'h00000cd0; 	    wdata_rom[  397] = 'hbad85d71; 	    wvalid_rom[  397] = 1; 
    i_addr_rom[  398] = 'h000000b8; 	    d_addr_rom[  398] = 'h00000f60; 	    wdata_rom[  398] = 'h293ddaca; 	    wvalid_rom[  398] = 0; 
    i_addr_rom[  399] = 'h000007a4; 	    d_addr_rom[  399] = 'h00000bfc; 	    wdata_rom[  399] = 'h6a85da8a; 	    wvalid_rom[  399] = 1; 
    i_addr_rom[  400] = 'h00000458; 	    d_addr_rom[  400] = 'h00000ab8; 	    wdata_rom[  400] = 'hb48ae587; 	    wvalid_rom[  400] = 0; 
    i_addr_rom[  401] = 'h00000784; 	    d_addr_rom[  401] = 'h00000ffc; 	    wdata_rom[  401] = 'ha69576ec; 	    wvalid_rom[  401] = 0; 
    i_addr_rom[  402] = 'h000004ac; 	    d_addr_rom[  402] = 'h00000a58; 	    wdata_rom[  402] = 'h149baeed; 	    wvalid_rom[  402] = 0; 
    i_addr_rom[  403] = 'h000007a8; 	    d_addr_rom[  403] = 'h000008ac; 	    wdata_rom[  403] = 'h7798c113; 	    wvalid_rom[  403] = 1; 
    i_addr_rom[  404] = 'h00000530; 	    d_addr_rom[  404] = 'h0000084c; 	    wdata_rom[  404] = 'h8d10ed0f; 	    wvalid_rom[  404] = 0; 
    i_addr_rom[  405] = 'h000003e4; 	    d_addr_rom[  405] = 'h00000c68; 	    wdata_rom[  405] = 'ha6a29d30; 	    wvalid_rom[  405] = 0; 
    i_addr_rom[  406] = 'h00000438; 	    d_addr_rom[  406] = 'h00000a20; 	    wdata_rom[  406] = 'hfbca29c8; 	    wvalid_rom[  406] = 0; 
    i_addr_rom[  407] = 'h000002cc; 	    d_addr_rom[  407] = 'h00000d08; 	    wdata_rom[  407] = 'h7ad8ca12; 	    wvalid_rom[  407] = 1; 
    i_addr_rom[  408] = 'h000001e8; 	    d_addr_rom[  408] = 'h00000bd0; 	    wdata_rom[  408] = 'ha09c7e32; 	    wvalid_rom[  408] = 1; 
    i_addr_rom[  409] = 'h000000b8; 	    d_addr_rom[  409] = 'h00000c2c; 	    wdata_rom[  409] = 'hae637550; 	    wvalid_rom[  409] = 1; 
    i_addr_rom[  410] = 'h000002ac; 	    d_addr_rom[  410] = 'h00000f9c; 	    wdata_rom[  410] = 'h8789ead0; 	    wvalid_rom[  410] = 0; 
    i_addr_rom[  411] = 'h00000378; 	    d_addr_rom[  411] = 'h0000084c; 	    wdata_rom[  411] = 'h5049032f; 	    wvalid_rom[  411] = 1; 
    i_addr_rom[  412] = 'h0000064c; 	    d_addr_rom[  412] = 'h00000ca8; 	    wdata_rom[  412] = 'hcc625d63; 	    wvalid_rom[  412] = 0; 
    i_addr_rom[  413] = 'h000001f8; 	    d_addr_rom[  413] = 'h00000fec; 	    wdata_rom[  413] = 'hb6e86c65; 	    wvalid_rom[  413] = 1; 
    i_addr_rom[  414] = 'h00000024; 	    d_addr_rom[  414] = 'h00000c94; 	    wdata_rom[  414] = 'h0e316aa2; 	    wvalid_rom[  414] = 0; 
    i_addr_rom[  415] = 'h000003f4; 	    d_addr_rom[  415] = 'h00000de4; 	    wdata_rom[  415] = 'hbfddbecc; 	    wvalid_rom[  415] = 1; 
    i_addr_rom[  416] = 'h000003a8; 	    d_addr_rom[  416] = 'h00000cc8; 	    wdata_rom[  416] = 'h2d1028a2; 	    wvalid_rom[  416] = 1; 
    i_addr_rom[  417] = 'h00000788; 	    d_addr_rom[  417] = 'h00000fd0; 	    wdata_rom[  417] = 'hc5e2b3a7; 	    wvalid_rom[  417] = 1; 
    i_addr_rom[  418] = 'h0000007c; 	    d_addr_rom[  418] = 'h00000e08; 	    wdata_rom[  418] = 'h3449e201; 	    wvalid_rom[  418] = 1; 
    i_addr_rom[  419] = 'h00000224; 	    d_addr_rom[  419] = 'h00000a44; 	    wdata_rom[  419] = 'h420d8a1a; 	    wvalid_rom[  419] = 1; 
    i_addr_rom[  420] = 'h00000764; 	    d_addr_rom[  420] = 'h00000ac8; 	    wdata_rom[  420] = 'hf0bbbc96; 	    wvalid_rom[  420] = 1; 
    i_addr_rom[  421] = 'h0000029c; 	    d_addr_rom[  421] = 'h00000e0c; 	    wdata_rom[  421] = 'h9ff3dd85; 	    wvalid_rom[  421] = 1; 
    i_addr_rom[  422] = 'h00000664; 	    d_addr_rom[  422] = 'h00000a44; 	    wdata_rom[  422] = 'headfedb5; 	    wvalid_rom[  422] = 1; 
    i_addr_rom[  423] = 'h0000040c; 	    d_addr_rom[  423] = 'h00000d04; 	    wdata_rom[  423] = 'hb547f0ae; 	    wvalid_rom[  423] = 0; 
    i_addr_rom[  424] = 'h00000354; 	    d_addr_rom[  424] = 'h00000898; 	    wdata_rom[  424] = 'hdfbfc56c; 	    wvalid_rom[  424] = 0; 
    i_addr_rom[  425] = 'h000001e0; 	    d_addr_rom[  425] = 'h00000f20; 	    wdata_rom[  425] = 'h78fe52a4; 	    wvalid_rom[  425] = 0; 
    i_addr_rom[  426] = 'h0000040c; 	    d_addr_rom[  426] = 'h00000fb0; 	    wdata_rom[  426] = 'h5d686d73; 	    wvalid_rom[  426] = 1; 
    i_addr_rom[  427] = 'h00000644; 	    d_addr_rom[  427] = 'h00000c30; 	    wdata_rom[  427] = 'hb650e22c; 	    wvalid_rom[  427] = 1; 
    i_addr_rom[  428] = 'h00000520; 	    d_addr_rom[  428] = 'h000008cc; 	    wdata_rom[  428] = 'heb69cb66; 	    wvalid_rom[  428] = 0; 
    i_addr_rom[  429] = 'h00000354; 	    d_addr_rom[  429] = 'h000009e0; 	    wdata_rom[  429] = 'h1f3d82b9; 	    wvalid_rom[  429] = 0; 
    i_addr_rom[  430] = 'h00000270; 	    d_addr_rom[  430] = 'h00000c08; 	    wdata_rom[  430] = 'hdf6c563b; 	    wvalid_rom[  430] = 1; 
    i_addr_rom[  431] = 'h00000784; 	    d_addr_rom[  431] = 'h000009e8; 	    wdata_rom[  431] = 'hf3a8a5c4; 	    wvalid_rom[  431] = 0; 
    i_addr_rom[  432] = 'h000002c8; 	    d_addr_rom[  432] = 'h0000089c; 	    wdata_rom[  432] = 'ha4853411; 	    wvalid_rom[  432] = 1; 
    i_addr_rom[  433] = 'h00000624; 	    d_addr_rom[  433] = 'h00000f84; 	    wdata_rom[  433] = 'h5a954b8d; 	    wvalid_rom[  433] = 0; 
    i_addr_rom[  434] = 'h00000370; 	    d_addr_rom[  434] = 'h00000f98; 	    wdata_rom[  434] = 'h1030311e; 	    wvalid_rom[  434] = 0; 
    i_addr_rom[  435] = 'h00000544; 	    d_addr_rom[  435] = 'h00000e58; 	    wdata_rom[  435] = 'h028ec881; 	    wvalid_rom[  435] = 0; 
    i_addr_rom[  436] = 'h00000164; 	    d_addr_rom[  436] = 'h00000af8; 	    wdata_rom[  436] = 'h91bb7520; 	    wvalid_rom[  436] = 1; 
    i_addr_rom[  437] = 'h00000198; 	    d_addr_rom[  437] = 'h00000d44; 	    wdata_rom[  437] = 'h6c557441; 	    wvalid_rom[  437] = 1; 
    i_addr_rom[  438] = 'h0000056c; 	    d_addr_rom[  438] = 'h000008f4; 	    wdata_rom[  438] = 'h09f24cd6; 	    wvalid_rom[  438] = 0; 
    i_addr_rom[  439] = 'h00000654; 	    d_addr_rom[  439] = 'h00000d50; 	    wdata_rom[  439] = 'h428c328e; 	    wvalid_rom[  439] = 1; 
    i_addr_rom[  440] = 'h00000664; 	    d_addr_rom[  440] = 'h00000958; 	    wdata_rom[  440] = 'h2bf013d2; 	    wvalid_rom[  440] = 0; 
    i_addr_rom[  441] = 'h0000062c; 	    d_addr_rom[  441] = 'h00000b94; 	    wdata_rom[  441] = 'hdf0966ba; 	    wvalid_rom[  441] = 1; 
    i_addr_rom[  442] = 'h00000178; 	    d_addr_rom[  442] = 'h00000a10; 	    wdata_rom[  442] = 'h531bbd32; 	    wvalid_rom[  442] = 1; 
    i_addr_rom[  443] = 'h00000130; 	    d_addr_rom[  443] = 'h00000af0; 	    wdata_rom[  443] = 'h3f601488; 	    wvalid_rom[  443] = 0; 
    i_addr_rom[  444] = 'h000003a8; 	    d_addr_rom[  444] = 'h00000a80; 	    wdata_rom[  444] = 'h7f811eb5; 	    wvalid_rom[  444] = 0; 
    i_addr_rom[  445] = 'h0000009c; 	    d_addr_rom[  445] = 'h00000cc4; 	    wdata_rom[  445] = 'h977db008; 	    wvalid_rom[  445] = 1; 
    i_addr_rom[  446] = 'h00000484; 	    d_addr_rom[  446] = 'h00000bbc; 	    wdata_rom[  446] = 'hb9121337; 	    wvalid_rom[  446] = 0; 
    i_addr_rom[  447] = 'h00000758; 	    d_addr_rom[  447] = 'h00000d18; 	    wdata_rom[  447] = 'h09398856; 	    wvalid_rom[  447] = 0; 
    i_addr_rom[  448] = 'h0000021c; 	    d_addr_rom[  448] = 'h00000cf8; 	    wdata_rom[  448] = 'h4c0b11e4; 	    wvalid_rom[  448] = 0; 
    i_addr_rom[  449] = 'h00000254; 	    d_addr_rom[  449] = 'h00000ab4; 	    wdata_rom[  449] = 'h90566e0e; 	    wvalid_rom[  449] = 0; 
    i_addr_rom[  450] = 'h00000374; 	    d_addr_rom[  450] = 'h00000b84; 	    wdata_rom[  450] = 'h1b85b2ce; 	    wvalid_rom[  450] = 1; 
    i_addr_rom[  451] = 'h00000308; 	    d_addr_rom[  451] = 'h00000e84; 	    wdata_rom[  451] = 'h181b7c8b; 	    wvalid_rom[  451] = 0; 
    i_addr_rom[  452] = 'h000007f8; 	    d_addr_rom[  452] = 'h0000098c; 	    wdata_rom[  452] = 'h66fc1667; 	    wvalid_rom[  452] = 0; 
    i_addr_rom[  453] = 'h00000444; 	    d_addr_rom[  453] = 'h00000a2c; 	    wdata_rom[  453] = 'h80859cc0; 	    wvalid_rom[  453] = 0; 
    i_addr_rom[  454] = 'h0000062c; 	    d_addr_rom[  454] = 'h00000f90; 	    wdata_rom[  454] = 'h026e5560; 	    wvalid_rom[  454] = 0; 
    i_addr_rom[  455] = 'h000006e0; 	    d_addr_rom[  455] = 'h00000f80; 	    wdata_rom[  455] = 'h87f6e3c2; 	    wvalid_rom[  455] = 1; 
    i_addr_rom[  456] = 'h00000704; 	    d_addr_rom[  456] = 'h00000ec4; 	    wdata_rom[  456] = 'h8d810e09; 	    wvalid_rom[  456] = 0; 
    i_addr_rom[  457] = 'h00000010; 	    d_addr_rom[  457] = 'h000008d0; 	    wdata_rom[  457] = 'h3dccdece; 	    wvalid_rom[  457] = 0; 
    i_addr_rom[  458] = 'h00000184; 	    d_addr_rom[  458] = 'h00000d90; 	    wdata_rom[  458] = 'h17438cf3; 	    wvalid_rom[  458] = 1; 
    i_addr_rom[  459] = 'h000004f8; 	    d_addr_rom[  459] = 'h00000ca8; 	    wdata_rom[  459] = 'h2da84190; 	    wvalid_rom[  459] = 1; 
    i_addr_rom[  460] = 'h000002b8; 	    d_addr_rom[  460] = 'h00000d34; 	    wdata_rom[  460] = 'h25927ff9; 	    wvalid_rom[  460] = 0; 
    i_addr_rom[  461] = 'h00000264; 	    d_addr_rom[  461] = 'h00000b50; 	    wdata_rom[  461] = 'h5f66d64e; 	    wvalid_rom[  461] = 1; 
    i_addr_rom[  462] = 'h000000d0; 	    d_addr_rom[  462] = 'h00000ad8; 	    wdata_rom[  462] = 'hff86c5ac; 	    wvalid_rom[  462] = 1; 
    i_addr_rom[  463] = 'h000002a8; 	    d_addr_rom[  463] = 'h000009a8; 	    wdata_rom[  463] = 'haa627519; 	    wvalid_rom[  463] = 0; 
    i_addr_rom[  464] = 'h00000040; 	    d_addr_rom[  464] = 'h00000bfc; 	    wdata_rom[  464] = 'hf28e4647; 	    wvalid_rom[  464] = 0; 
    i_addr_rom[  465] = 'h00000044; 	    d_addr_rom[  465] = 'h00000f90; 	    wdata_rom[  465] = 'hf9669b0c; 	    wvalid_rom[  465] = 1; 
    i_addr_rom[  466] = 'h00000460; 	    d_addr_rom[  466] = 'h00000908; 	    wdata_rom[  466] = 'h38c69993; 	    wvalid_rom[  466] = 1; 
    i_addr_rom[  467] = 'h00000118; 	    d_addr_rom[  467] = 'h00000cdc; 	    wdata_rom[  467] = 'hfb93b505; 	    wvalid_rom[  467] = 0; 
    i_addr_rom[  468] = 'h000002fc; 	    d_addr_rom[  468] = 'h00000b08; 	    wdata_rom[  468] = 'hefc2d866; 	    wvalid_rom[  468] = 1; 
    i_addr_rom[  469] = 'h00000740; 	    d_addr_rom[  469] = 'h00000c58; 	    wdata_rom[  469] = 'h713b033f; 	    wvalid_rom[  469] = 1; 
    i_addr_rom[  470] = 'h00000760; 	    d_addr_rom[  470] = 'h000008a8; 	    wdata_rom[  470] = 'hbc58af03; 	    wvalid_rom[  470] = 0; 
    i_addr_rom[  471] = 'h00000438; 	    d_addr_rom[  471] = 'h00000aa8; 	    wdata_rom[  471] = 'hed78f115; 	    wvalid_rom[  471] = 0; 
    i_addr_rom[  472] = 'h000001ec; 	    d_addr_rom[  472] = 'h00000e28; 	    wdata_rom[  472] = 'hb48d830a; 	    wvalid_rom[  472] = 0; 
    i_addr_rom[  473] = 'h000006fc; 	    d_addr_rom[  473] = 'h00000db8; 	    wdata_rom[  473] = 'h5bd278f4; 	    wvalid_rom[  473] = 1; 
    i_addr_rom[  474] = 'h00000778; 	    d_addr_rom[  474] = 'h00000dac; 	    wdata_rom[  474] = 'hd0b67fa7; 	    wvalid_rom[  474] = 1; 
    i_addr_rom[  475] = 'h000004e4; 	    d_addr_rom[  475] = 'h00000cf0; 	    wdata_rom[  475] = 'h9ea53452; 	    wvalid_rom[  475] = 0; 
    i_addr_rom[  476] = 'h000003cc; 	    d_addr_rom[  476] = 'h00000860; 	    wdata_rom[  476] = 'h24ff2301; 	    wvalid_rom[  476] = 0; 
    i_addr_rom[  477] = 'h00000664; 	    d_addr_rom[  477] = 'h00000ef4; 	    wdata_rom[  477] = 'he910d9b1; 	    wvalid_rom[  477] = 0; 
    i_addr_rom[  478] = 'h00000588; 	    d_addr_rom[  478] = 'h000008dc; 	    wdata_rom[  478] = 'h158989e3; 	    wvalid_rom[  478] = 1; 
    i_addr_rom[  479] = 'h00000228; 	    d_addr_rom[  479] = 'h00000bac; 	    wdata_rom[  479] = 'hffd9fb73; 	    wvalid_rom[  479] = 1; 
    i_addr_rom[  480] = 'h0000073c; 	    d_addr_rom[  480] = 'h00000fa8; 	    wdata_rom[  480] = 'he55a05d2; 	    wvalid_rom[  480] = 0; 
    i_addr_rom[  481] = 'h0000043c; 	    d_addr_rom[  481] = 'h00000d54; 	    wdata_rom[  481] = 'hfb6b32e8; 	    wvalid_rom[  481] = 0; 
    i_addr_rom[  482] = 'h000000bc; 	    d_addr_rom[  482] = 'h00000bf8; 	    wdata_rom[  482] = 'he15671d6; 	    wvalid_rom[  482] = 1; 
    i_addr_rom[  483] = 'h000005a0; 	    d_addr_rom[  483] = 'h00000aec; 	    wdata_rom[  483] = 'h9a482bb3; 	    wvalid_rom[  483] = 0; 
    i_addr_rom[  484] = 'h00000504; 	    d_addr_rom[  484] = 'h00000fec; 	    wdata_rom[  484] = 'hffe32893; 	    wvalid_rom[  484] = 1; 
    i_addr_rom[  485] = 'h0000056c; 	    d_addr_rom[  485] = 'h00000b34; 	    wdata_rom[  485] = 'h820d2fbd; 	    wvalid_rom[  485] = 1; 
    i_addr_rom[  486] = 'h00000778; 	    d_addr_rom[  486] = 'h00000bb4; 	    wdata_rom[  486] = 'hb6399155; 	    wvalid_rom[  486] = 0; 
    i_addr_rom[  487] = 'h00000140; 	    d_addr_rom[  487] = 'h00000bac; 	    wdata_rom[  487] = 'h035ee8da; 	    wvalid_rom[  487] = 0; 
    i_addr_rom[  488] = 'h00000188; 	    d_addr_rom[  488] = 'h00000d94; 	    wdata_rom[  488] = 'hd0a2a72a; 	    wvalid_rom[  488] = 1; 
    i_addr_rom[  489] = 'h00000750; 	    d_addr_rom[  489] = 'h00000f14; 	    wdata_rom[  489] = 'he7da207d; 	    wvalid_rom[  489] = 1; 
    i_addr_rom[  490] = 'h00000708; 	    d_addr_rom[  490] = 'h0000085c; 	    wdata_rom[  490] = 'hfed3d6a2; 	    wvalid_rom[  490] = 0; 
    i_addr_rom[  491] = 'h000002d4; 	    d_addr_rom[  491] = 'h00000bec; 	    wdata_rom[  491] = 'h53b89727; 	    wvalid_rom[  491] = 0; 
    i_addr_rom[  492] = 'h000003d0; 	    d_addr_rom[  492] = 'h00000a10; 	    wdata_rom[  492] = 'h33d90b8f; 	    wvalid_rom[  492] = 1; 
    i_addr_rom[  493] = 'h00000670; 	    d_addr_rom[  493] = 'h0000085c; 	    wdata_rom[  493] = 'h09fa6fda; 	    wvalid_rom[  493] = 1; 
    i_addr_rom[  494] = 'h000005d0; 	    d_addr_rom[  494] = 'h00000c18; 	    wdata_rom[  494] = 'ha1adc72e; 	    wvalid_rom[  494] = 0; 
    i_addr_rom[  495] = 'h000004f4; 	    d_addr_rom[  495] = 'h00000984; 	    wdata_rom[  495] = 'h697f62d7; 	    wvalid_rom[  495] = 1; 
    i_addr_rom[  496] = 'h0000032c; 	    d_addr_rom[  496] = 'h000009f8; 	    wdata_rom[  496] = 'h34ac56fa; 	    wvalid_rom[  496] = 0; 
    i_addr_rom[  497] = 'h00000284; 	    d_addr_rom[  497] = 'h00000e84; 	    wdata_rom[  497] = 'h9a523096; 	    wvalid_rom[  497] = 0; 
    i_addr_rom[  498] = 'h00000180; 	    d_addr_rom[  498] = 'h00000b50; 	    wdata_rom[  498] = 'h8d946578; 	    wvalid_rom[  498] = 1; 
    i_addr_rom[  499] = 'h000000b4; 	    d_addr_rom[  499] = 'h00000bf8; 	    wdata_rom[  499] = 'h1317ea7c; 	    wvalid_rom[  499] = 1; 
    i_addr_rom[  500] = 'h00000614; 	    d_addr_rom[  500] = 'h00000e5c; 	    wdata_rom[  500] = 'h812ab067; 	    wvalid_rom[  500] = 1; 
    i_addr_rom[  501] = 'h0000020c; 	    d_addr_rom[  501] = 'h00000d58; 	    wdata_rom[  501] = 'h67ee1d94; 	    wvalid_rom[  501] = 0; 
    i_addr_rom[  502] = 'h00000428; 	    d_addr_rom[  502] = 'h00000b94; 	    wdata_rom[  502] = 'h42ec8963; 	    wvalid_rom[  502] = 1; 
    i_addr_rom[  503] = 'h000000d0; 	    d_addr_rom[  503] = 'h000008a4; 	    wdata_rom[  503] = 'ha85bc37e; 	    wvalid_rom[  503] = 1; 
    i_addr_rom[  504] = 'h00000088; 	    d_addr_rom[  504] = 'h00000cfc; 	    wdata_rom[  504] = 'h981395e4; 	    wvalid_rom[  504] = 1; 
    i_addr_rom[  505] = 'h00000460; 	    d_addr_rom[  505] = 'h00000fb8; 	    wdata_rom[  505] = 'h0c818285; 	    wvalid_rom[  505] = 1; 
    i_addr_rom[  506] = 'h000005dc; 	    d_addr_rom[  506] = 'h00000f18; 	    wdata_rom[  506] = 'hf55b94f3; 	    wvalid_rom[  506] = 0; 
    i_addr_rom[  507] = 'h00000764; 	    d_addr_rom[  507] = 'h00000d30; 	    wdata_rom[  507] = 'h01c80ed4; 	    wvalid_rom[  507] = 0; 
    i_addr_rom[  508] = 'h00000274; 	    d_addr_rom[  508] = 'h00000a90; 	    wdata_rom[  508] = 'h72290f48; 	    wvalid_rom[  508] = 1; 
    i_addr_rom[  509] = 'h00000064; 	    d_addr_rom[  509] = 'h00000da0; 	    wdata_rom[  509] = 'he00cc83f; 	    wvalid_rom[  509] = 0; 
    i_addr_rom[  510] = 'h000007b4; 	    d_addr_rom[  510] = 'h00000f98; 	    wdata_rom[  510] = 'h29a10b17; 	    wvalid_rom[  510] = 0; 
    i_addr_rom[  511] = 'h000003a8; 	    d_addr_rom[  511] = 'h000009cc; 	    wdata_rom[  511] = 'h1aabac7a; 	    wvalid_rom[  511] = 0; 
    i_addr_rom[  512] = 'h00000268; 	    d_addr_rom[  512] = 'h00000be0; 	    wdata_rom[  512] = 'h7edccdaa; 	    wvalid_rom[  512] = 1; 
    i_addr_rom[  513] = 'h00000214; 	    d_addr_rom[  513] = 'h00000d7c; 	    wdata_rom[  513] = 'h4538bfaa; 	    wvalid_rom[  513] = 0; 
    i_addr_rom[  514] = 'h000007c0; 	    d_addr_rom[  514] = 'h00000e20; 	    wdata_rom[  514] = 'h5d392e2c; 	    wvalid_rom[  514] = 1; 
    i_addr_rom[  515] = 'h00000714; 	    d_addr_rom[  515] = 'h00000ce0; 	    wdata_rom[  515] = 'ha7c764df; 	    wvalid_rom[  515] = 0; 
    i_addr_rom[  516] = 'h00000450; 	    d_addr_rom[  516] = 'h00000884; 	    wdata_rom[  516] = 'h3dc31f85; 	    wvalid_rom[  516] = 0; 
    i_addr_rom[  517] = 'h000000f0; 	    d_addr_rom[  517] = 'h000009ac; 	    wdata_rom[  517] = 'h29512b60; 	    wvalid_rom[  517] = 1; 
    i_addr_rom[  518] = 'h0000057c; 	    d_addr_rom[  518] = 'h00000d6c; 	    wdata_rom[  518] = 'h2d67e00a; 	    wvalid_rom[  518] = 0; 
    i_addr_rom[  519] = 'h000006b8; 	    d_addr_rom[  519] = 'h00000e30; 	    wdata_rom[  519] = 'h0f7d4567; 	    wvalid_rom[  519] = 1; 
    i_addr_rom[  520] = 'h000003d0; 	    d_addr_rom[  520] = 'h00000e0c; 	    wdata_rom[  520] = 'hb9022c37; 	    wvalid_rom[  520] = 0; 
    i_addr_rom[  521] = 'h00000334; 	    d_addr_rom[  521] = 'h00000990; 	    wdata_rom[  521] = 'hf0221124; 	    wvalid_rom[  521] = 1; 
    i_addr_rom[  522] = 'h00000318; 	    d_addr_rom[  522] = 'h00000e4c; 	    wdata_rom[  522] = 'h27427cb1; 	    wvalid_rom[  522] = 0; 
    i_addr_rom[  523] = 'h000005a0; 	    d_addr_rom[  523] = 'h00000f00; 	    wdata_rom[  523] = 'h18309efe; 	    wvalid_rom[  523] = 0; 
    i_addr_rom[  524] = 'h00000124; 	    d_addr_rom[  524] = 'h00000cac; 	    wdata_rom[  524] = 'hf0c54ca8; 	    wvalid_rom[  524] = 1; 
    i_addr_rom[  525] = 'h0000072c; 	    d_addr_rom[  525] = 'h00000e98; 	    wdata_rom[  525] = 'h3133e4fc; 	    wvalid_rom[  525] = 1; 
    i_addr_rom[  526] = 'h00000688; 	    d_addr_rom[  526] = 'h00000eac; 	    wdata_rom[  526] = 'hb7166164; 	    wvalid_rom[  526] = 0; 
    i_addr_rom[  527] = 'h000001cc; 	    d_addr_rom[  527] = 'h0000094c; 	    wdata_rom[  527] = 'h534e0da3; 	    wvalid_rom[  527] = 1; 
    i_addr_rom[  528] = 'h00000724; 	    d_addr_rom[  528] = 'h00000de0; 	    wdata_rom[  528] = 'h425d896c; 	    wvalid_rom[  528] = 1; 
    i_addr_rom[  529] = 'h00000178; 	    d_addr_rom[  529] = 'h00000ab0; 	    wdata_rom[  529] = 'h16f55126; 	    wvalid_rom[  529] = 0; 
    i_addr_rom[  530] = 'h00000398; 	    d_addr_rom[  530] = 'h00000be0; 	    wdata_rom[  530] = 'hbd271bce; 	    wvalid_rom[  530] = 0; 
    i_addr_rom[  531] = 'h00000300; 	    d_addr_rom[  531] = 'h00000acc; 	    wdata_rom[  531] = 'hf09d51d2; 	    wvalid_rom[  531] = 0; 
    i_addr_rom[  532] = 'h00000100; 	    d_addr_rom[  532] = 'h000008ec; 	    wdata_rom[  532] = 'h9428b210; 	    wvalid_rom[  532] = 0; 
    i_addr_rom[  533] = 'h00000478; 	    d_addr_rom[  533] = 'h00000914; 	    wdata_rom[  533] = 'hdef28428; 	    wvalid_rom[  533] = 1; 
    i_addr_rom[  534] = 'h0000079c; 	    d_addr_rom[  534] = 'h00000ec8; 	    wdata_rom[  534] = 'hf1d5c830; 	    wvalid_rom[  534] = 0; 
    i_addr_rom[  535] = 'h0000066c; 	    d_addr_rom[  535] = 'h00000970; 	    wdata_rom[  535] = 'h6bfffaca; 	    wvalid_rom[  535] = 1; 
    i_addr_rom[  536] = 'h00000074; 	    d_addr_rom[  536] = 'h00000f84; 	    wdata_rom[  536] = 'h0cc966ef; 	    wvalid_rom[  536] = 1; 
    i_addr_rom[  537] = 'h00000070; 	    d_addr_rom[  537] = 'h00000c0c; 	    wdata_rom[  537] = 'h2c543ad7; 	    wvalid_rom[  537] = 1; 
    i_addr_rom[  538] = 'h000007f4; 	    d_addr_rom[  538] = 'h00000e00; 	    wdata_rom[  538] = 'h608c2321; 	    wvalid_rom[  538] = 1; 
    i_addr_rom[  539] = 'h0000078c; 	    d_addr_rom[  539] = 'h00000f90; 	    wdata_rom[  539] = 'h1cc69b03; 	    wvalid_rom[  539] = 1; 
    i_addr_rom[  540] = 'h000005c8; 	    d_addr_rom[  540] = 'h00000d50; 	    wdata_rom[  540] = 'h65434740; 	    wvalid_rom[  540] = 0; 
    i_addr_rom[  541] = 'h00000110; 	    d_addr_rom[  541] = 'h00000b54; 	    wdata_rom[  541] = 'h1f2252d4; 	    wvalid_rom[  541] = 0; 
    i_addr_rom[  542] = 'h000007cc; 	    d_addr_rom[  542] = 'h00000a28; 	    wdata_rom[  542] = 'h3b4e1922; 	    wvalid_rom[  542] = 1; 
    i_addr_rom[  543] = 'h000003bc; 	    d_addr_rom[  543] = 'h00000ee4; 	    wdata_rom[  543] = 'h52208a87; 	    wvalid_rom[  543] = 1; 
    i_addr_rom[  544] = 'h00000284; 	    d_addr_rom[  544] = 'h000009f4; 	    wdata_rom[  544] = 'h3f67c070; 	    wvalid_rom[  544] = 1; 
    i_addr_rom[  545] = 'h000001b8; 	    d_addr_rom[  545] = 'h0000099c; 	    wdata_rom[  545] = 'h14e7ce1a; 	    wvalid_rom[  545] = 0; 
    i_addr_rom[  546] = 'h000001d8; 	    d_addr_rom[  546] = 'h000008f0; 	    wdata_rom[  546] = 'h42df15c7; 	    wvalid_rom[  546] = 0; 
    i_addr_rom[  547] = 'h00000424; 	    d_addr_rom[  547] = 'h000008b4; 	    wdata_rom[  547] = 'h73442252; 	    wvalid_rom[  547] = 0; 
    i_addr_rom[  548] = 'h000005f8; 	    d_addr_rom[  548] = 'h00000924; 	    wdata_rom[  548] = 'he04d36b2; 	    wvalid_rom[  548] = 0; 
    i_addr_rom[  549] = 'h000003fc; 	    d_addr_rom[  549] = 'h00000d14; 	    wdata_rom[  549] = 'h4bb9bf94; 	    wvalid_rom[  549] = 0; 
    i_addr_rom[  550] = 'h00000248; 	    d_addr_rom[  550] = 'h00000870; 	    wdata_rom[  550] = 'h9b26459c; 	    wvalid_rom[  550] = 1; 
    i_addr_rom[  551] = 'h00000000; 	    d_addr_rom[  551] = 'h00000b58; 	    wdata_rom[  551] = 'h9786d06a; 	    wvalid_rom[  551] = 0; 
    i_addr_rom[  552] = 'h00000060; 	    d_addr_rom[  552] = 'h00000ffc; 	    wdata_rom[  552] = 'hae4654db; 	    wvalid_rom[  552] = 1; 
    i_addr_rom[  553] = 'h00000618; 	    d_addr_rom[  553] = 'h00000890; 	    wdata_rom[  553] = 'h640237d6; 	    wvalid_rom[  553] = 1; 
    i_addr_rom[  554] = 'h000006fc; 	    d_addr_rom[  554] = 'h00000cbc; 	    wdata_rom[  554] = 'h16b02ca1; 	    wvalid_rom[  554] = 1; 
    i_addr_rom[  555] = 'h00000108; 	    d_addr_rom[  555] = 'h0000095c; 	    wdata_rom[  555] = 'h327fd13a; 	    wvalid_rom[  555] = 1; 
    i_addr_rom[  556] = 'h0000068c; 	    d_addr_rom[  556] = 'h00000e48; 	    wdata_rom[  556] = 'h402f83fa; 	    wvalid_rom[  556] = 1; 
    i_addr_rom[  557] = 'h00000200; 	    d_addr_rom[  557] = 'h00000c6c; 	    wdata_rom[  557] = 'h9a5bb6cc; 	    wvalid_rom[  557] = 0; 
    i_addr_rom[  558] = 'h00000018; 	    d_addr_rom[  558] = 'h00000838; 	    wdata_rom[  558] = 'he31d8254; 	    wvalid_rom[  558] = 1; 
    i_addr_rom[  559] = 'h000004b0; 	    d_addr_rom[  559] = 'h00000934; 	    wdata_rom[  559] = 'h29310ee2; 	    wvalid_rom[  559] = 1; 
    i_addr_rom[  560] = 'h00000220; 	    d_addr_rom[  560] = 'h00000818; 	    wdata_rom[  560] = 'h27eb7e21; 	    wvalid_rom[  560] = 0; 
    i_addr_rom[  561] = 'h00000600; 	    d_addr_rom[  561] = 'h00000b2c; 	    wdata_rom[  561] = 'h57660399; 	    wvalid_rom[  561] = 0; 
    i_addr_rom[  562] = 'h000004dc; 	    d_addr_rom[  562] = 'h00000e48; 	    wdata_rom[  562] = 'h151323b1; 	    wvalid_rom[  562] = 1; 
    i_addr_rom[  563] = 'h00000298; 	    d_addr_rom[  563] = 'h00000d04; 	    wdata_rom[  563] = 'h1700c46e; 	    wvalid_rom[  563] = 1; 
    i_addr_rom[  564] = 'h000007c8; 	    d_addr_rom[  564] = 'h00000de8; 	    wdata_rom[  564] = 'hd477ad90; 	    wvalid_rom[  564] = 1; 
    i_addr_rom[  565] = 'h00000630; 	    d_addr_rom[  565] = 'h00000d60; 	    wdata_rom[  565] = 'h06c08fe9; 	    wvalid_rom[  565] = 1; 
    i_addr_rom[  566] = 'h000005d8; 	    d_addr_rom[  566] = 'h00000c48; 	    wdata_rom[  566] = 'hbd877a16; 	    wvalid_rom[  566] = 0; 
    i_addr_rom[  567] = 'h0000070c; 	    d_addr_rom[  567] = 'h00000f90; 	    wdata_rom[  567] = 'he84c6e6a; 	    wvalid_rom[  567] = 1; 
    i_addr_rom[  568] = 'h00000470; 	    d_addr_rom[  568] = 'h00000b0c; 	    wdata_rom[  568] = 'h36a7c62d; 	    wvalid_rom[  568] = 0; 
    i_addr_rom[  569] = 'h000003f4; 	    d_addr_rom[  569] = 'h00000d98; 	    wdata_rom[  569] = 'h66898690; 	    wvalid_rom[  569] = 0; 
    i_addr_rom[  570] = 'h000005a8; 	    d_addr_rom[  570] = 'h00000b38; 	    wdata_rom[  570] = 'h17e30da8; 	    wvalid_rom[  570] = 1; 
    i_addr_rom[  571] = 'h00000168; 	    d_addr_rom[  571] = 'h00000818; 	    wdata_rom[  571] = 'h793bce8d; 	    wvalid_rom[  571] = 1; 
    i_addr_rom[  572] = 'h0000042c; 	    d_addr_rom[  572] = 'h00000eb0; 	    wdata_rom[  572] = 'h04698ecf; 	    wvalid_rom[  572] = 1; 
    i_addr_rom[  573] = 'h0000079c; 	    d_addr_rom[  573] = 'h00000bc0; 	    wdata_rom[  573] = 'h5d29fae5; 	    wvalid_rom[  573] = 0; 
    i_addr_rom[  574] = 'h000004c0; 	    d_addr_rom[  574] = 'h00000d48; 	    wdata_rom[  574] = 'h485fe35e; 	    wvalid_rom[  574] = 0; 
    i_addr_rom[  575] = 'h00000104; 	    d_addr_rom[  575] = 'h0000083c; 	    wdata_rom[  575] = 'he686d7b0; 	    wvalid_rom[  575] = 1; 
    i_addr_rom[  576] = 'h000006a4; 	    d_addr_rom[  576] = 'h00000d08; 	    wdata_rom[  576] = 'hb08ed809; 	    wvalid_rom[  576] = 1; 
    i_addr_rom[  577] = 'h0000079c; 	    d_addr_rom[  577] = 'h00000be8; 	    wdata_rom[  577] = 'hc8068926; 	    wvalid_rom[  577] = 0; 
    i_addr_rom[  578] = 'h00000114; 	    d_addr_rom[  578] = 'h00000a38; 	    wdata_rom[  578] = 'hc3b6258d; 	    wvalid_rom[  578] = 0; 
    i_addr_rom[  579] = 'h00000698; 	    d_addr_rom[  579] = 'h00000c34; 	    wdata_rom[  579] = 'h25a5e068; 	    wvalid_rom[  579] = 1; 
    i_addr_rom[  580] = 'h000005b4; 	    d_addr_rom[  580] = 'h00000da4; 	    wdata_rom[  580] = 'hf5b08712; 	    wvalid_rom[  580] = 1; 
    i_addr_rom[  581] = 'h0000004c; 	    d_addr_rom[  581] = 'h00000bc0; 	    wdata_rom[  581] = 'he92ab92d; 	    wvalid_rom[  581] = 1; 
    i_addr_rom[  582] = 'h00000050; 	    d_addr_rom[  582] = 'h000008e4; 	    wdata_rom[  582] = 'h55bf8226; 	    wvalid_rom[  582] = 1; 
    i_addr_rom[  583] = 'h00000788; 	    d_addr_rom[  583] = 'h00000eec; 	    wdata_rom[  583] = 'h337761d7; 	    wvalid_rom[  583] = 0; 
    i_addr_rom[  584] = 'h000004f8; 	    d_addr_rom[  584] = 'h00000ddc; 	    wdata_rom[  584] = 'h532ee801; 	    wvalid_rom[  584] = 1; 
    i_addr_rom[  585] = 'h000006e4; 	    d_addr_rom[  585] = 'h00000cc8; 	    wdata_rom[  585] = 'hd895234e; 	    wvalid_rom[  585] = 1; 
    i_addr_rom[  586] = 'h000001b8; 	    d_addr_rom[  586] = 'h00000d50; 	    wdata_rom[  586] = 'h1757a726; 	    wvalid_rom[  586] = 1; 
    i_addr_rom[  587] = 'h000001f8; 	    d_addr_rom[  587] = 'h00000940; 	    wdata_rom[  587] = 'h1b7a8122; 	    wvalid_rom[  587] = 1; 
    i_addr_rom[  588] = 'h00000108; 	    d_addr_rom[  588] = 'h00000e5c; 	    wdata_rom[  588] = 'h7d53d658; 	    wvalid_rom[  588] = 1; 
    i_addr_rom[  589] = 'h00000244; 	    d_addr_rom[  589] = 'h00000f58; 	    wdata_rom[  589] = 'h1b8f5567; 	    wvalid_rom[  589] = 1; 
    i_addr_rom[  590] = 'h00000378; 	    d_addr_rom[  590] = 'h00000f90; 	    wdata_rom[  590] = 'h228b755b; 	    wvalid_rom[  590] = 1; 
    i_addr_rom[  591] = 'h00000594; 	    d_addr_rom[  591] = 'h00000954; 	    wdata_rom[  591] = 'h32d1a259; 	    wvalid_rom[  591] = 1; 
    i_addr_rom[  592] = 'h000006cc; 	    d_addr_rom[  592] = 'h00000a64; 	    wdata_rom[  592] = 'h25e509b6; 	    wvalid_rom[  592] = 0; 
    i_addr_rom[  593] = 'h00000280; 	    d_addr_rom[  593] = 'h00000d58; 	    wdata_rom[  593] = 'he4df3bea; 	    wvalid_rom[  593] = 0; 
    i_addr_rom[  594] = 'h000006ac; 	    d_addr_rom[  594] = 'h00000920; 	    wdata_rom[  594] = 'h886717fe; 	    wvalid_rom[  594] = 0; 
    i_addr_rom[  595] = 'h0000062c; 	    d_addr_rom[  595] = 'h00000ecc; 	    wdata_rom[  595] = 'h3d905a45; 	    wvalid_rom[  595] = 0; 
    i_addr_rom[  596] = 'h00000628; 	    d_addr_rom[  596] = 'h00000bec; 	    wdata_rom[  596] = 'h4ec98a2c; 	    wvalid_rom[  596] = 0; 
    i_addr_rom[  597] = 'h000003c8; 	    d_addr_rom[  597] = 'h00000a6c; 	    wdata_rom[  597] = 'he0672fa3; 	    wvalid_rom[  597] = 1; 
    i_addr_rom[  598] = 'h0000048c; 	    d_addr_rom[  598] = 'h00000f38; 	    wdata_rom[  598] = 'h8cc510f2; 	    wvalid_rom[  598] = 1; 
    i_addr_rom[  599] = 'h0000030c; 	    d_addr_rom[  599] = 'h00000e10; 	    wdata_rom[  599] = 'hf8c59fcb; 	    wvalid_rom[  599] = 1; 
    i_addr_rom[  600] = 'h00000424; 	    d_addr_rom[  600] = 'h00000ee4; 	    wdata_rom[  600] = 'h76cc5df0; 	    wvalid_rom[  600] = 1; 
    i_addr_rom[  601] = 'h00000254; 	    d_addr_rom[  601] = 'h00000b1c; 	    wdata_rom[  601] = 'h70c3e74c; 	    wvalid_rom[  601] = 0; 
    i_addr_rom[  602] = 'h00000498; 	    d_addr_rom[  602] = 'h00000868; 	    wdata_rom[  602] = 'h68694d55; 	    wvalid_rom[  602] = 0; 
    i_addr_rom[  603] = 'h00000078; 	    d_addr_rom[  603] = 'h00000c08; 	    wdata_rom[  603] = 'hda2e7367; 	    wvalid_rom[  603] = 0; 
    i_addr_rom[  604] = 'h00000324; 	    d_addr_rom[  604] = 'h000009b8; 	    wdata_rom[  604] = 'h7237b75e; 	    wvalid_rom[  604] = 0; 
    i_addr_rom[  605] = 'h00000510; 	    d_addr_rom[  605] = 'h00000e2c; 	    wdata_rom[  605] = 'h47dc6499; 	    wvalid_rom[  605] = 1; 
    i_addr_rom[  606] = 'h000003f0; 	    d_addr_rom[  606] = 'h00000d74; 	    wdata_rom[  606] = 'h0b17005a; 	    wvalid_rom[  606] = 1; 
    i_addr_rom[  607] = 'h00000524; 	    d_addr_rom[  607] = 'h00000af4; 	    wdata_rom[  607] = 'h41e8b385; 	    wvalid_rom[  607] = 1; 
    i_addr_rom[  608] = 'h00000050; 	    d_addr_rom[  608] = 'h00000b10; 	    wdata_rom[  608] = 'h49966e5b; 	    wvalid_rom[  608] = 1; 
    i_addr_rom[  609] = 'h00000328; 	    d_addr_rom[  609] = 'h0000092c; 	    wdata_rom[  609] = 'h9dbac375; 	    wvalid_rom[  609] = 0; 
    i_addr_rom[  610] = 'h00000474; 	    d_addr_rom[  610] = 'h00000f10; 	    wdata_rom[  610] = 'ha034a441; 	    wvalid_rom[  610] = 0; 
    i_addr_rom[  611] = 'h000002f0; 	    d_addr_rom[  611] = 'h000009d0; 	    wdata_rom[  611] = 'h27b49997; 	    wvalid_rom[  611] = 0; 
    i_addr_rom[  612] = 'h000003a4; 	    d_addr_rom[  612] = 'h00000818; 	    wdata_rom[  612] = 'h4d7f3eaa; 	    wvalid_rom[  612] = 1; 
    i_addr_rom[  613] = 'h0000050c; 	    d_addr_rom[  613] = 'h00000eac; 	    wdata_rom[  613] = 'h90d37e0d; 	    wvalid_rom[  613] = 1; 
    i_addr_rom[  614] = 'h00000604; 	    d_addr_rom[  614] = 'h00000b38; 	    wdata_rom[  614] = 'h8b24ca4a; 	    wvalid_rom[  614] = 1; 
    i_addr_rom[  615] = 'h000003cc; 	    d_addr_rom[  615] = 'h00000e64; 	    wdata_rom[  615] = 'h4f74744f; 	    wvalid_rom[  615] = 1; 
    i_addr_rom[  616] = 'h000006f8; 	    d_addr_rom[  616] = 'h000008a4; 	    wdata_rom[  616] = 'h5baca976; 	    wvalid_rom[  616] = 1; 
    i_addr_rom[  617] = 'h0000078c; 	    d_addr_rom[  617] = 'h00000cac; 	    wdata_rom[  617] = 'h7ecaec2c; 	    wvalid_rom[  617] = 1; 
    i_addr_rom[  618] = 'h00000164; 	    d_addr_rom[  618] = 'h00000d14; 	    wdata_rom[  618] = 'h650fc1e6; 	    wvalid_rom[  618] = 1; 
    i_addr_rom[  619] = 'h00000054; 	    d_addr_rom[  619] = 'h00000ca8; 	    wdata_rom[  619] = 'h82ad5136; 	    wvalid_rom[  619] = 0; 
    i_addr_rom[  620] = 'h000000e0; 	    d_addr_rom[  620] = 'h00000f30; 	    wdata_rom[  620] = 'hbab6d089; 	    wvalid_rom[  620] = 0; 
    i_addr_rom[  621] = 'h000002f0; 	    d_addr_rom[  621] = 'h00000860; 	    wdata_rom[  621] = 'ha2b37278; 	    wvalid_rom[  621] = 0; 
    i_addr_rom[  622] = 'h00000530; 	    d_addr_rom[  622] = 'h00000da0; 	    wdata_rom[  622] = 'h172b6a0c; 	    wvalid_rom[  622] = 1; 
    i_addr_rom[  623] = 'h000006ec; 	    d_addr_rom[  623] = 'h00000eac; 	    wdata_rom[  623] = 'hefecc3f7; 	    wvalid_rom[  623] = 1; 
    i_addr_rom[  624] = 'h00000750; 	    d_addr_rom[  624] = 'h00000e44; 	    wdata_rom[  624] = 'h52f41d7c; 	    wvalid_rom[  624] = 1; 
    i_addr_rom[  625] = 'h000002c8; 	    d_addr_rom[  625] = 'h000009e0; 	    wdata_rom[  625] = 'h58d9c3b0; 	    wvalid_rom[  625] = 0; 
    i_addr_rom[  626] = 'h0000025c; 	    d_addr_rom[  626] = 'h00000d80; 	    wdata_rom[  626] = 'h139e6951; 	    wvalid_rom[  626] = 0; 
    i_addr_rom[  627] = 'h0000026c; 	    d_addr_rom[  627] = 'h00000fbc; 	    wdata_rom[  627] = 'hdde54f7a; 	    wvalid_rom[  627] = 1; 
    i_addr_rom[  628] = 'h000005dc; 	    d_addr_rom[  628] = 'h00000fb0; 	    wdata_rom[  628] = 'hef8dc06e; 	    wvalid_rom[  628] = 1; 
    i_addr_rom[  629] = 'h0000052c; 	    d_addr_rom[  629] = 'h000008c0; 	    wdata_rom[  629] = 'h4bbc526f; 	    wvalid_rom[  629] = 0; 
    i_addr_rom[  630] = 'h000001b0; 	    d_addr_rom[  630] = 'h00000f9c; 	    wdata_rom[  630] = 'h683ceade; 	    wvalid_rom[  630] = 1; 
    i_addr_rom[  631] = 'h000003b4; 	    d_addr_rom[  631] = 'h000008fc; 	    wdata_rom[  631] = 'hf8ec07b1; 	    wvalid_rom[  631] = 0; 
    i_addr_rom[  632] = 'h000001d8; 	    d_addr_rom[  632] = 'h00000a40; 	    wdata_rom[  632] = 'ha99b68c1; 	    wvalid_rom[  632] = 1; 
    i_addr_rom[  633] = 'h0000077c; 	    d_addr_rom[  633] = 'h00000d94; 	    wdata_rom[  633] = 'hd9ca4f91; 	    wvalid_rom[  633] = 1; 
    i_addr_rom[  634] = 'h0000054c; 	    d_addr_rom[  634] = 'h00000b90; 	    wdata_rom[  634] = 'h9767d451; 	    wvalid_rom[  634] = 0; 
    i_addr_rom[  635] = 'h000007bc; 	    d_addr_rom[  635] = 'h00000eac; 	    wdata_rom[  635] = 'h7cf59939; 	    wvalid_rom[  635] = 1; 
    i_addr_rom[  636] = 'h00000204; 	    d_addr_rom[  636] = 'h0000098c; 	    wdata_rom[  636] = 'hd625dbeb; 	    wvalid_rom[  636] = 1; 
    i_addr_rom[  637] = 'h0000068c; 	    d_addr_rom[  637] = 'h00000ab8; 	    wdata_rom[  637] = 'h4e01a177; 	    wvalid_rom[  637] = 0; 
    i_addr_rom[  638] = 'h00000668; 	    d_addr_rom[  638] = 'h00000af0; 	    wdata_rom[  638] = 'h61703896; 	    wvalid_rom[  638] = 0; 
    i_addr_rom[  639] = 'h00000244; 	    d_addr_rom[  639] = 'h00000b90; 	    wdata_rom[  639] = 'hf045e9d5; 	    wvalid_rom[  639] = 1; 
    i_addr_rom[  640] = 'h00000630; 	    d_addr_rom[  640] = 'h00000ab4; 	    wdata_rom[  640] = 'h79ad7b6d; 	    wvalid_rom[  640] = 0; 
    i_addr_rom[  641] = 'h00000488; 	    d_addr_rom[  641] = 'h00000f38; 	    wdata_rom[  641] = 'h8825df86; 	    wvalid_rom[  641] = 0; 
    i_addr_rom[  642] = 'h00000314; 	    d_addr_rom[  642] = 'h00000920; 	    wdata_rom[  642] = 'h3ae64b99; 	    wvalid_rom[  642] = 0; 
    i_addr_rom[  643] = 'h000005d0; 	    d_addr_rom[  643] = 'h00000c90; 	    wdata_rom[  643] = 'h60f41064; 	    wvalid_rom[  643] = 1; 
    i_addr_rom[  644] = 'h0000024c; 	    d_addr_rom[  644] = 'h00000e24; 	    wdata_rom[  644] = 'h666b4ae3; 	    wvalid_rom[  644] = 0; 
    i_addr_rom[  645] = 'h000005d8; 	    d_addr_rom[  645] = 'h00000b90; 	    wdata_rom[  645] = 'h52866278; 	    wvalid_rom[  645] = 0; 
    i_addr_rom[  646] = 'h00000308; 	    d_addr_rom[  646] = 'h00000ed8; 	    wdata_rom[  646] = 'hc9fb4518; 	    wvalid_rom[  646] = 1; 
    i_addr_rom[  647] = 'h000005f0; 	    d_addr_rom[  647] = 'h00000cc4; 	    wdata_rom[  647] = 'h1d8afcef; 	    wvalid_rom[  647] = 1; 
    i_addr_rom[  648] = 'h000006c4; 	    d_addr_rom[  648] = 'h0000088c; 	    wdata_rom[  648] = 'h06d562cb; 	    wvalid_rom[  648] = 1; 
    i_addr_rom[  649] = 'h0000005c; 	    d_addr_rom[  649] = 'h00000eec; 	    wdata_rom[  649] = 'h2658b586; 	    wvalid_rom[  649] = 1; 
    i_addr_rom[  650] = 'h00000348; 	    d_addr_rom[  650] = 'h00000c2c; 	    wdata_rom[  650] = 'h325c0a33; 	    wvalid_rom[  650] = 0; 
    i_addr_rom[  651] = 'h000006bc; 	    d_addr_rom[  651] = 'h000008b4; 	    wdata_rom[  651] = 'h33ab2aff; 	    wvalid_rom[  651] = 1; 
    i_addr_rom[  652] = 'h00000200; 	    d_addr_rom[  652] = 'h00000f34; 	    wdata_rom[  652] = 'h83f68877; 	    wvalid_rom[  652] = 1; 
    i_addr_rom[  653] = 'h00000100; 	    d_addr_rom[  653] = 'h00000bd0; 	    wdata_rom[  653] = 'h7e820463; 	    wvalid_rom[  653] = 0; 
    i_addr_rom[  654] = 'h000007b8; 	    d_addr_rom[  654] = 'h00000ef8; 	    wdata_rom[  654] = 'h82e88d83; 	    wvalid_rom[  654] = 1; 
    i_addr_rom[  655] = 'h00000780; 	    d_addr_rom[  655] = 'h00000d78; 	    wdata_rom[  655] = 'hb62a911a; 	    wvalid_rom[  655] = 0; 
    i_addr_rom[  656] = 'h00000138; 	    d_addr_rom[  656] = 'h00000d78; 	    wdata_rom[  656] = 'hecd9704b; 	    wvalid_rom[  656] = 0; 
    i_addr_rom[  657] = 'h000004a0; 	    d_addr_rom[  657] = 'h00000bf4; 	    wdata_rom[  657] = 'h6cc199f8; 	    wvalid_rom[  657] = 0; 
    i_addr_rom[  658] = 'h000006d4; 	    d_addr_rom[  658] = 'h00000d08; 	    wdata_rom[  658] = 'heb3588d6; 	    wvalid_rom[  658] = 1; 
    i_addr_rom[  659] = 'h00000110; 	    d_addr_rom[  659] = 'h00000b08; 	    wdata_rom[  659] = 'h175d5452; 	    wvalid_rom[  659] = 0; 
    i_addr_rom[  660] = 'h000000e0; 	    d_addr_rom[  660] = 'h00000bb0; 	    wdata_rom[  660] = 'h9b9da915; 	    wvalid_rom[  660] = 0; 
    i_addr_rom[  661] = 'h00000528; 	    d_addr_rom[  661] = 'h00000c08; 	    wdata_rom[  661] = 'h1d7b3983; 	    wvalid_rom[  661] = 0; 
    i_addr_rom[  662] = 'h000002b4; 	    d_addr_rom[  662] = 'h00000a8c; 	    wdata_rom[  662] = 'haa8a8f3a; 	    wvalid_rom[  662] = 0; 
    i_addr_rom[  663] = 'h000000c0; 	    d_addr_rom[  663] = 'h00000dcc; 	    wdata_rom[  663] = 'h5c7e2d5c; 	    wvalid_rom[  663] = 0; 
    i_addr_rom[  664] = 'h00000314; 	    d_addr_rom[  664] = 'h00000848; 	    wdata_rom[  664] = 'h30c721ee; 	    wvalid_rom[  664] = 1; 
    i_addr_rom[  665] = 'h00000220; 	    d_addr_rom[  665] = 'h00000f0c; 	    wdata_rom[  665] = 'h32edc64f; 	    wvalid_rom[  665] = 0; 
    i_addr_rom[  666] = 'h00000098; 	    d_addr_rom[  666] = 'h00000874; 	    wdata_rom[  666] = 'h786d94ee; 	    wvalid_rom[  666] = 1; 
    i_addr_rom[  667] = 'h00000644; 	    d_addr_rom[  667] = 'h00000ff8; 	    wdata_rom[  667] = 'hf2287561; 	    wvalid_rom[  667] = 1; 
    i_addr_rom[  668] = 'h000006d0; 	    d_addr_rom[  668] = 'h00000e7c; 	    wdata_rom[  668] = 'h53434847; 	    wvalid_rom[  668] = 0; 
    i_addr_rom[  669] = 'h000004d8; 	    d_addr_rom[  669] = 'h00000af0; 	    wdata_rom[  669] = 'h1db2764d; 	    wvalid_rom[  669] = 0; 
    i_addr_rom[  670] = 'h000005b0; 	    d_addr_rom[  670] = 'h000008c4; 	    wdata_rom[  670] = 'h4c4cd1f5; 	    wvalid_rom[  670] = 0; 
    i_addr_rom[  671] = 'h0000046c; 	    d_addr_rom[  671] = 'h00000cc8; 	    wdata_rom[  671] = 'ha4020fd6; 	    wvalid_rom[  671] = 0; 
    i_addr_rom[  672] = 'h0000035c; 	    d_addr_rom[  672] = 'h00000e48; 	    wdata_rom[  672] = 'hd0202f09; 	    wvalid_rom[  672] = 1; 
    i_addr_rom[  673] = 'h0000025c; 	    d_addr_rom[  673] = 'h00000ba8; 	    wdata_rom[  673] = 'h831eef2a; 	    wvalid_rom[  673] = 1; 
    i_addr_rom[  674] = 'h0000063c; 	    d_addr_rom[  674] = 'h00000bbc; 	    wdata_rom[  674] = 'h160b16a3; 	    wvalid_rom[  674] = 1; 
    i_addr_rom[  675] = 'h000007f0; 	    d_addr_rom[  675] = 'h00000dd8; 	    wdata_rom[  675] = 'h718f97b9; 	    wvalid_rom[  675] = 1; 
    i_addr_rom[  676] = 'h00000458; 	    d_addr_rom[  676] = 'h00000910; 	    wdata_rom[  676] = 'h6ce5a1f3; 	    wvalid_rom[  676] = 1; 
    i_addr_rom[  677] = 'h000001b0; 	    d_addr_rom[  677] = 'h0000099c; 	    wdata_rom[  677] = 'h4bbce149; 	    wvalid_rom[  677] = 0; 
    i_addr_rom[  678] = 'h000004c0; 	    d_addr_rom[  678] = 'h00000eb0; 	    wdata_rom[  678] = 'h1be17111; 	    wvalid_rom[  678] = 1; 
    i_addr_rom[  679] = 'h0000001c; 	    d_addr_rom[  679] = 'h00000ec4; 	    wdata_rom[  679] = 'hd8b1024c; 	    wvalid_rom[  679] = 0; 
    i_addr_rom[  680] = 'h0000049c; 	    d_addr_rom[  680] = 'h00000b98; 	    wdata_rom[  680] = 'h98d4a29b; 	    wvalid_rom[  680] = 0; 
    i_addr_rom[  681] = 'h0000029c; 	    d_addr_rom[  681] = 'h00000ab8; 	    wdata_rom[  681] = 'hcd321223; 	    wvalid_rom[  681] = 1; 
    i_addr_rom[  682] = 'h00000008; 	    d_addr_rom[  682] = 'h00000c70; 	    wdata_rom[  682] = 'h23431ece; 	    wvalid_rom[  682] = 1; 
    i_addr_rom[  683] = 'h000000c4; 	    d_addr_rom[  683] = 'h00000ab8; 	    wdata_rom[  683] = 'h329ce4f4; 	    wvalid_rom[  683] = 1; 
    i_addr_rom[  684] = 'h000002dc; 	    d_addr_rom[  684] = 'h00000cf8; 	    wdata_rom[  684] = 'h398c5446; 	    wvalid_rom[  684] = 1; 
    i_addr_rom[  685] = 'h00000048; 	    d_addr_rom[  685] = 'h00000ed8; 	    wdata_rom[  685] = 'h6ed2d6be; 	    wvalid_rom[  685] = 0; 
    i_addr_rom[  686] = 'h00000490; 	    d_addr_rom[  686] = 'h00000d78; 	    wdata_rom[  686] = 'h9fe3629e; 	    wvalid_rom[  686] = 1; 
    i_addr_rom[  687] = 'h00000500; 	    d_addr_rom[  687] = 'h000008e4; 	    wdata_rom[  687] = 'h80e49049; 	    wvalid_rom[  687] = 1; 
    i_addr_rom[  688] = 'h00000780; 	    d_addr_rom[  688] = 'h0000086c; 	    wdata_rom[  688] = 'h8d189a2c; 	    wvalid_rom[  688] = 1; 
    i_addr_rom[  689] = 'h00000144; 	    d_addr_rom[  689] = 'h00000c0c; 	    wdata_rom[  689] = 'h0ab94ae9; 	    wvalid_rom[  689] = 1; 
    i_addr_rom[  690] = 'h000002d0; 	    d_addr_rom[  690] = 'h0000096c; 	    wdata_rom[  690] = 'h7e14d8b8; 	    wvalid_rom[  690] = 1; 
    i_addr_rom[  691] = 'h00000664; 	    d_addr_rom[  691] = 'h00000e20; 	    wdata_rom[  691] = 'h75d436e5; 	    wvalid_rom[  691] = 0; 
    i_addr_rom[  692] = 'h000002b4; 	    d_addr_rom[  692] = 'h00000f10; 	    wdata_rom[  692] = 'h20355448; 	    wvalid_rom[  692] = 0; 
    i_addr_rom[  693] = 'h000000e0; 	    d_addr_rom[  693] = 'h0000081c; 	    wdata_rom[  693] = 'h2824ce88; 	    wvalid_rom[  693] = 1; 
    i_addr_rom[  694] = 'h00000470; 	    d_addr_rom[  694] = 'h00000d98; 	    wdata_rom[  694] = 'h340c5be8; 	    wvalid_rom[  694] = 1; 
    i_addr_rom[  695] = 'h00000250; 	    d_addr_rom[  695] = 'h00000afc; 	    wdata_rom[  695] = 'h88f7a66e; 	    wvalid_rom[  695] = 1; 
    i_addr_rom[  696] = 'h000007e8; 	    d_addr_rom[  696] = 'h00000bcc; 	    wdata_rom[  696] = 'h198ed70e; 	    wvalid_rom[  696] = 0; 
    i_addr_rom[  697] = 'h00000298; 	    d_addr_rom[  697] = 'h00000c0c; 	    wdata_rom[  697] = 'h19ab7b8a; 	    wvalid_rom[  697] = 0; 
    i_addr_rom[  698] = 'h0000040c; 	    d_addr_rom[  698] = 'h00000ca4; 	    wdata_rom[  698] = 'hfb51d441; 	    wvalid_rom[  698] = 0; 
    i_addr_rom[  699] = 'h00000664; 	    d_addr_rom[  699] = 'h00000940; 	    wdata_rom[  699] = 'hcef1a4cb; 	    wvalid_rom[  699] = 1; 
    i_addr_rom[  700] = 'h00000210; 	    d_addr_rom[  700] = 'h000008d4; 	    wdata_rom[  700] = 'hc2100f66; 	    wvalid_rom[  700] = 1; 
    i_addr_rom[  701] = 'h000003c4; 	    d_addr_rom[  701] = 'h000009e0; 	    wdata_rom[  701] = 'hd6569082; 	    wvalid_rom[  701] = 1; 
    i_addr_rom[  702] = 'h000002b8; 	    d_addr_rom[  702] = 'h00000c4c; 	    wdata_rom[  702] = 'h56f15ab3; 	    wvalid_rom[  702] = 0; 
    i_addr_rom[  703] = 'h00000720; 	    d_addr_rom[  703] = 'h00000ec4; 	    wdata_rom[  703] = 'he9e7320e; 	    wvalid_rom[  703] = 1; 
    i_addr_rom[  704] = 'h00000390; 	    d_addr_rom[  704] = 'h00000b7c; 	    wdata_rom[  704] = 'h103d7c3e; 	    wvalid_rom[  704] = 1; 
    i_addr_rom[  705] = 'h0000031c; 	    d_addr_rom[  705] = 'h000008a8; 	    wdata_rom[  705] = 'he7bb40ad; 	    wvalid_rom[  705] = 1; 
    i_addr_rom[  706] = 'h000005f8; 	    d_addr_rom[  706] = 'h00000fe0; 	    wdata_rom[  706] = 'hfdc56d9a; 	    wvalid_rom[  706] = 1; 
    i_addr_rom[  707] = 'h00000008; 	    d_addr_rom[  707] = 'h00000f64; 	    wdata_rom[  707] = 'h2d62a90c; 	    wvalid_rom[  707] = 0; 
    i_addr_rom[  708] = 'h000004c4; 	    d_addr_rom[  708] = 'h00000aa8; 	    wdata_rom[  708] = 'h079a95de; 	    wvalid_rom[  708] = 0; 
    i_addr_rom[  709] = 'h00000304; 	    d_addr_rom[  709] = 'h00000c00; 	    wdata_rom[  709] = 'hb9d8b1f3; 	    wvalid_rom[  709] = 0; 
    i_addr_rom[  710] = 'h0000043c; 	    d_addr_rom[  710] = 'h00000d7c; 	    wdata_rom[  710] = 'h67c05981; 	    wvalid_rom[  710] = 0; 
    i_addr_rom[  711] = 'h0000026c; 	    d_addr_rom[  711] = 'h00000fcc; 	    wdata_rom[  711] = 'ha2398fd8; 	    wvalid_rom[  711] = 0; 
    i_addr_rom[  712] = 'h000006d0; 	    d_addr_rom[  712] = 'h00000998; 	    wdata_rom[  712] = 'hac871e78; 	    wvalid_rom[  712] = 0; 
    i_addr_rom[  713] = 'h0000019c; 	    d_addr_rom[  713] = 'h000009ec; 	    wdata_rom[  713] = 'h01bcaeda; 	    wvalid_rom[  713] = 0; 
    i_addr_rom[  714] = 'h000005d0; 	    d_addr_rom[  714] = 'h00000e34; 	    wdata_rom[  714] = 'he68c321e; 	    wvalid_rom[  714] = 1; 
    i_addr_rom[  715] = 'h000006b0; 	    d_addr_rom[  715] = 'h00000f90; 	    wdata_rom[  715] = 'he3cb5574; 	    wvalid_rom[  715] = 1; 
    i_addr_rom[  716] = 'h00000354; 	    d_addr_rom[  716] = 'h000008b4; 	    wdata_rom[  716] = 'h48ca2b17; 	    wvalid_rom[  716] = 0; 
    i_addr_rom[  717] = 'h00000524; 	    d_addr_rom[  717] = 'h00000cf4; 	    wdata_rom[  717] = 'hc7badab9; 	    wvalid_rom[  717] = 1; 
    i_addr_rom[  718] = 'h00000758; 	    d_addr_rom[  718] = 'h00000978; 	    wdata_rom[  718] = 'hdbeafc0a; 	    wvalid_rom[  718] = 1; 
    i_addr_rom[  719] = 'h00000328; 	    d_addr_rom[  719] = 'h00000f68; 	    wdata_rom[  719] = 'h299d6bba; 	    wvalid_rom[  719] = 1; 
    i_addr_rom[  720] = 'h00000628; 	    d_addr_rom[  720] = 'h00000978; 	    wdata_rom[  720] = 'h836d4b61; 	    wvalid_rom[  720] = 1; 
    i_addr_rom[  721] = 'h00000000; 	    d_addr_rom[  721] = 'h00000868; 	    wdata_rom[  721] = 'hc57f4f0a; 	    wvalid_rom[  721] = 0; 
    i_addr_rom[  722] = 'h000007e8; 	    d_addr_rom[  722] = 'h00000f34; 	    wdata_rom[  722] = 'hafec4179; 	    wvalid_rom[  722] = 0; 
    i_addr_rom[  723] = 'h0000009c; 	    d_addr_rom[  723] = 'h00000b28; 	    wdata_rom[  723] = 'he4845b73; 	    wvalid_rom[  723] = 0; 
    i_addr_rom[  724] = 'h000000f0; 	    d_addr_rom[  724] = 'h00000920; 	    wdata_rom[  724] = 'h6590c243; 	    wvalid_rom[  724] = 1; 
    i_addr_rom[  725] = 'h00000720; 	    d_addr_rom[  725] = 'h00000904; 	    wdata_rom[  725] = 'h2dc4c59b; 	    wvalid_rom[  725] = 0; 
    i_addr_rom[  726] = 'h000007a4; 	    d_addr_rom[  726] = 'h00000ba4; 	    wdata_rom[  726] = 'h7368b4c3; 	    wvalid_rom[  726] = 1; 
    i_addr_rom[  727] = 'h000006c0; 	    d_addr_rom[  727] = 'h00000eb0; 	    wdata_rom[  727] = 'ha9d454f3; 	    wvalid_rom[  727] = 1; 
    i_addr_rom[  728] = 'h000006b0; 	    d_addr_rom[  728] = 'h00000c10; 	    wdata_rom[  728] = 'h7d9e4dbd; 	    wvalid_rom[  728] = 0; 
    i_addr_rom[  729] = 'h00000694; 	    d_addr_rom[  729] = 'h00000b28; 	    wdata_rom[  729] = 'hcd25d576; 	    wvalid_rom[  729] = 0; 
    i_addr_rom[  730] = 'h000004a0; 	    d_addr_rom[  730] = 'h000009cc; 	    wdata_rom[  730] = 'hea5aca7d; 	    wvalid_rom[  730] = 1; 
    i_addr_rom[  731] = 'h000000a4; 	    d_addr_rom[  731] = 'h00000964; 	    wdata_rom[  731] = 'hd01daf9d; 	    wvalid_rom[  731] = 1; 
    i_addr_rom[  732] = 'h00000280; 	    d_addr_rom[  732] = 'h00000c40; 	    wdata_rom[  732] = 'h49bc14a6; 	    wvalid_rom[  732] = 0; 
    i_addr_rom[  733] = 'h000001c8; 	    d_addr_rom[  733] = 'h000009d8; 	    wdata_rom[  733] = 'h28012281; 	    wvalid_rom[  733] = 0; 
    i_addr_rom[  734] = 'h0000071c; 	    d_addr_rom[  734] = 'h00000c58; 	    wdata_rom[  734] = 'hd7cf9ac7; 	    wvalid_rom[  734] = 0; 
    i_addr_rom[  735] = 'h00000768; 	    d_addr_rom[  735] = 'h00000c00; 	    wdata_rom[  735] = 'hec1a8ad8; 	    wvalid_rom[  735] = 1; 
    i_addr_rom[  736] = 'h000004ec; 	    d_addr_rom[  736] = 'h00000ca4; 	    wdata_rom[  736] = 'hab8177f3; 	    wvalid_rom[  736] = 1; 
    i_addr_rom[  737] = 'h00000064; 	    d_addr_rom[  737] = 'h00000904; 	    wdata_rom[  737] = 'h2a1feb3e; 	    wvalid_rom[  737] = 1; 
    i_addr_rom[  738] = 'h000007b8; 	    d_addr_rom[  738] = 'h00000bb4; 	    wdata_rom[  738] = 'h7ee23670; 	    wvalid_rom[  738] = 1; 
    i_addr_rom[  739] = 'h0000020c; 	    d_addr_rom[  739] = 'h00000f30; 	    wdata_rom[  739] = 'h1ca24ac2; 	    wvalid_rom[  739] = 0; 
    i_addr_rom[  740] = 'h000007e4; 	    d_addr_rom[  740] = 'h00000c04; 	    wdata_rom[  740] = 'hbc0f7f70; 	    wvalid_rom[  740] = 0; 
    i_addr_rom[  741] = 'h00000418; 	    d_addr_rom[  741] = 'h00000df8; 	    wdata_rom[  741] = 'h3c6b45d4; 	    wvalid_rom[  741] = 1; 
    i_addr_rom[  742] = 'h00000344; 	    d_addr_rom[  742] = 'h00000b84; 	    wdata_rom[  742] = 'h92dcd436; 	    wvalid_rom[  742] = 0; 
    i_addr_rom[  743] = 'h00000664; 	    d_addr_rom[  743] = 'h00000e2c; 	    wdata_rom[  743] = 'h3cec4e40; 	    wvalid_rom[  743] = 0; 
    i_addr_rom[  744] = 'h0000050c; 	    d_addr_rom[  744] = 'h00000fcc; 	    wdata_rom[  744] = 'h04827284; 	    wvalid_rom[  744] = 0; 
    i_addr_rom[  745] = 'h0000008c; 	    d_addr_rom[  745] = 'h00000e24; 	    wdata_rom[  745] = 'h0d595df2; 	    wvalid_rom[  745] = 0; 
    i_addr_rom[  746] = 'h000007bc; 	    d_addr_rom[  746] = 'h00000c18; 	    wdata_rom[  746] = 'h9c4e4a34; 	    wvalid_rom[  746] = 0; 
    i_addr_rom[  747] = 'h000002a0; 	    d_addr_rom[  747] = 'h00000fc8; 	    wdata_rom[  747] = 'h6c21a1b6; 	    wvalid_rom[  747] = 0; 
    i_addr_rom[  748] = 'h00000394; 	    d_addr_rom[  748] = 'h00000cfc; 	    wdata_rom[  748] = 'h5df49eec; 	    wvalid_rom[  748] = 0; 
    i_addr_rom[  749] = 'h000002e8; 	    d_addr_rom[  749] = 'h00000888; 	    wdata_rom[  749] = 'hc297ab81; 	    wvalid_rom[  749] = 1; 
    i_addr_rom[  750] = 'h00000018; 	    d_addr_rom[  750] = 'h00000b68; 	    wdata_rom[  750] = 'h228e95c6; 	    wvalid_rom[  750] = 1; 
    i_addr_rom[  751] = 'h0000004c; 	    d_addr_rom[  751] = 'h00000b24; 	    wdata_rom[  751] = 'hf279ed3a; 	    wvalid_rom[  751] = 1; 
    i_addr_rom[  752] = 'h000006f4; 	    d_addr_rom[  752] = 'h00000a40; 	    wdata_rom[  752] = 'haccdc3c0; 	    wvalid_rom[  752] = 0; 
    i_addr_rom[  753] = 'h0000001c; 	    d_addr_rom[  753] = 'h00000c0c; 	    wdata_rom[  753] = 'hb577245b; 	    wvalid_rom[  753] = 0; 
    i_addr_rom[  754] = 'h00000048; 	    d_addr_rom[  754] = 'h00000e50; 	    wdata_rom[  754] = 'he41d72c8; 	    wvalid_rom[  754] = 1; 
    i_addr_rom[  755] = 'h0000018c; 	    d_addr_rom[  755] = 'h00000974; 	    wdata_rom[  755] = 'h6ab1250c; 	    wvalid_rom[  755] = 0; 
    i_addr_rom[  756] = 'h00000328; 	    d_addr_rom[  756] = 'h00000e38; 	    wdata_rom[  756] = 'hecfe184b; 	    wvalid_rom[  756] = 0; 
    i_addr_rom[  757] = 'h00000388; 	    d_addr_rom[  757] = 'h00000c54; 	    wdata_rom[  757] = 'h28fc7ef5; 	    wvalid_rom[  757] = 0; 
    i_addr_rom[  758] = 'h0000040c; 	    d_addr_rom[  758] = 'h00000e7c; 	    wdata_rom[  758] = 'h56ac4217; 	    wvalid_rom[  758] = 1; 
    i_addr_rom[  759] = 'h00000578; 	    d_addr_rom[  759] = 'h00000fa0; 	    wdata_rom[  759] = 'h56e75fe0; 	    wvalid_rom[  759] = 0; 
    i_addr_rom[  760] = 'h0000019c; 	    d_addr_rom[  760] = 'h00000e74; 	    wdata_rom[  760] = 'hf6688089; 	    wvalid_rom[  760] = 0; 
    i_addr_rom[  761] = 'h000004ac; 	    d_addr_rom[  761] = 'h00000d4c; 	    wdata_rom[  761] = 'h0a24cc3f; 	    wvalid_rom[  761] = 1; 
    i_addr_rom[  762] = 'h00000270; 	    d_addr_rom[  762] = 'h0000095c; 	    wdata_rom[  762] = 'h70ec1f0e; 	    wvalid_rom[  762] = 1; 
    i_addr_rom[  763] = 'h000002dc; 	    d_addr_rom[  763] = 'h00000edc; 	    wdata_rom[  763] = 'h92ecd089; 	    wvalid_rom[  763] = 0; 
    i_addr_rom[  764] = 'h00000498; 	    d_addr_rom[  764] = 'h00000ad0; 	    wdata_rom[  764] = 'h13569df8; 	    wvalid_rom[  764] = 1; 
    i_addr_rom[  765] = 'h000003b8; 	    d_addr_rom[  765] = 'h00000b20; 	    wdata_rom[  765] = 'hf9753fed; 	    wvalid_rom[  765] = 1; 
    i_addr_rom[  766] = 'h000005a8; 	    d_addr_rom[  766] = 'h00000d70; 	    wdata_rom[  766] = 'h8695cc26; 	    wvalid_rom[  766] = 1; 
    i_addr_rom[  767] = 'h000005c0; 	    d_addr_rom[  767] = 'h00000a90; 	    wdata_rom[  767] = 'heee6dd96; 	    wvalid_rom[  767] = 0; 
    i_addr_rom[  768] = 'h000004e4; 	    d_addr_rom[  768] = 'h00000de8; 	    wdata_rom[  768] = 'h2eed9d7e; 	    wvalid_rom[  768] = 1; 
    i_addr_rom[  769] = 'h000007e0; 	    d_addr_rom[  769] = 'h000008fc; 	    wdata_rom[  769] = 'h8e4d8427; 	    wvalid_rom[  769] = 1; 
    i_addr_rom[  770] = 'h00000364; 	    d_addr_rom[  770] = 'h00000c00; 	    wdata_rom[  770] = 'h988b68d8; 	    wvalid_rom[  770] = 0; 
    i_addr_rom[  771] = 'h00000388; 	    d_addr_rom[  771] = 'h00000ea0; 	    wdata_rom[  771] = 'h4870b16b; 	    wvalid_rom[  771] = 0; 
    i_addr_rom[  772] = 'h00000144; 	    d_addr_rom[  772] = 'h00000854; 	    wdata_rom[  772] = 'hcd823a79; 	    wvalid_rom[  772] = 0; 
    i_addr_rom[  773] = 'h000006e8; 	    d_addr_rom[  773] = 'h00000c34; 	    wdata_rom[  773] = 'hb90765d6; 	    wvalid_rom[  773] = 1; 
    i_addr_rom[  774] = 'h000002d4; 	    d_addr_rom[  774] = 'h00000ce0; 	    wdata_rom[  774] = 'h39da9c25; 	    wvalid_rom[  774] = 0; 
    i_addr_rom[  775] = 'h000002f4; 	    d_addr_rom[  775] = 'h00000fd4; 	    wdata_rom[  775] = 'h901dd650; 	    wvalid_rom[  775] = 1; 
    i_addr_rom[  776] = 'h00000260; 	    d_addr_rom[  776] = 'h0000099c; 	    wdata_rom[  776] = 'h5d6f94bc; 	    wvalid_rom[  776] = 1; 
    i_addr_rom[  777] = 'h000002b0; 	    d_addr_rom[  777] = 'h00000c6c; 	    wdata_rom[  777] = 'h96642d3b; 	    wvalid_rom[  777] = 1; 
    i_addr_rom[  778] = 'h0000030c; 	    d_addr_rom[  778] = 'h0000092c; 	    wdata_rom[  778] = 'h1ff03d4d; 	    wvalid_rom[  778] = 0; 
    i_addr_rom[  779] = 'h000006f0; 	    d_addr_rom[  779] = 'h00000fc8; 	    wdata_rom[  779] = 'h0c623aaf; 	    wvalid_rom[  779] = 0; 
    i_addr_rom[  780] = 'h00000320; 	    d_addr_rom[  780] = 'h00000bf8; 	    wdata_rom[  780] = 'h9d700eeb; 	    wvalid_rom[  780] = 1; 
    i_addr_rom[  781] = 'h000000e0; 	    d_addr_rom[  781] = 'h00000cb0; 	    wdata_rom[  781] = 'h500dd987; 	    wvalid_rom[  781] = 1; 
    i_addr_rom[  782] = 'h0000021c; 	    d_addr_rom[  782] = 'h00000c38; 	    wdata_rom[  782] = 'h013d015d; 	    wvalid_rom[  782] = 0; 
    i_addr_rom[  783] = 'h000001ec; 	    d_addr_rom[  783] = 'h00000bc8; 	    wdata_rom[  783] = 'hcf6f7679; 	    wvalid_rom[  783] = 0; 
    i_addr_rom[  784] = 'h000002dc; 	    d_addr_rom[  784] = 'h0000096c; 	    wdata_rom[  784] = 'had6baf04; 	    wvalid_rom[  784] = 0; 
    i_addr_rom[  785] = 'h0000063c; 	    d_addr_rom[  785] = 'h00000d0c; 	    wdata_rom[  785] = 'hbb36972d; 	    wvalid_rom[  785] = 1; 
    i_addr_rom[  786] = 'h00000144; 	    d_addr_rom[  786] = 'h00000e78; 	    wdata_rom[  786] = 'hf41976b2; 	    wvalid_rom[  786] = 0; 
    i_addr_rom[  787] = 'h00000038; 	    d_addr_rom[  787] = 'h00000ce0; 	    wdata_rom[  787] = 'h0999ed3c; 	    wvalid_rom[  787] = 1; 
    i_addr_rom[  788] = 'h00000208; 	    d_addr_rom[  788] = 'h00000c98; 	    wdata_rom[  788] = 'h3a3d6c6b; 	    wvalid_rom[  788] = 1; 
    i_addr_rom[  789] = 'h0000062c; 	    d_addr_rom[  789] = 'h00000cf4; 	    wdata_rom[  789] = 'h203cbd89; 	    wvalid_rom[  789] = 1; 
    i_addr_rom[  790] = 'h00000690; 	    d_addr_rom[  790] = 'h00000894; 	    wdata_rom[  790] = 'h35d2473c; 	    wvalid_rom[  790] = 1; 
    i_addr_rom[  791] = 'h000004a8; 	    d_addr_rom[  791] = 'h000008b0; 	    wdata_rom[  791] = 'he1c7901b; 	    wvalid_rom[  791] = 1; 
    i_addr_rom[  792] = 'h000003f4; 	    d_addr_rom[  792] = 'h000008bc; 	    wdata_rom[  792] = 'h80db5013; 	    wvalid_rom[  792] = 0; 
    i_addr_rom[  793] = 'h000003d4; 	    d_addr_rom[  793] = 'h00000a64; 	    wdata_rom[  793] = 'h6f831bf3; 	    wvalid_rom[  793] = 1; 
    i_addr_rom[  794] = 'h000002bc; 	    d_addr_rom[  794] = 'h00000a38; 	    wdata_rom[  794] = 'h92c58890; 	    wvalid_rom[  794] = 1; 
    i_addr_rom[  795] = 'h00000798; 	    d_addr_rom[  795] = 'h00000870; 	    wdata_rom[  795] = 'hba862dac; 	    wvalid_rom[  795] = 1; 
    i_addr_rom[  796] = 'h00000030; 	    d_addr_rom[  796] = 'h00000aa8; 	    wdata_rom[  796] = 'h8a6dfd62; 	    wvalid_rom[  796] = 1; 
    i_addr_rom[  797] = 'h000005a8; 	    d_addr_rom[  797] = 'h00000938; 	    wdata_rom[  797] = 'h05a86b8b; 	    wvalid_rom[  797] = 1; 
    i_addr_rom[  798] = 'h000005c8; 	    d_addr_rom[  798] = 'h00000c28; 	    wdata_rom[  798] = 'h2eda7f37; 	    wvalid_rom[  798] = 0; 
    i_addr_rom[  799] = 'h00000604; 	    d_addr_rom[  799] = 'h00000984; 	    wdata_rom[  799] = 'h242893ed; 	    wvalid_rom[  799] = 0; 
    i_addr_rom[  800] = 'h00000184; 	    d_addr_rom[  800] = 'h00000a08; 	    wdata_rom[  800] = 'h4cb95a4f; 	    wvalid_rom[  800] = 0; 
    i_addr_rom[  801] = 'h000006b4; 	    d_addr_rom[  801] = 'h00000ab8; 	    wdata_rom[  801] = 'h58642322; 	    wvalid_rom[  801] = 0; 
    i_addr_rom[  802] = 'h000001a0; 	    d_addr_rom[  802] = 'h00000da8; 	    wdata_rom[  802] = 'h2a2166a5; 	    wvalid_rom[  802] = 1; 
    i_addr_rom[  803] = 'h0000008c; 	    d_addr_rom[  803] = 'h00000c8c; 	    wdata_rom[  803] = 'h0ebd7b4b; 	    wvalid_rom[  803] = 1; 
    i_addr_rom[  804] = 'h00000438; 	    d_addr_rom[  804] = 'h00000c8c; 	    wdata_rom[  804] = 'hfe508ae7; 	    wvalid_rom[  804] = 0; 
    i_addr_rom[  805] = 'h000001b8; 	    d_addr_rom[  805] = 'h00000c40; 	    wdata_rom[  805] = 'hb6fc63bf; 	    wvalid_rom[  805] = 1; 
    i_addr_rom[  806] = 'h000006ac; 	    d_addr_rom[  806] = 'h00000e48; 	    wdata_rom[  806] = 'h94141b3c; 	    wvalid_rom[  806] = 0; 
    i_addr_rom[  807] = 'h0000073c; 	    d_addr_rom[  807] = 'h00000a34; 	    wdata_rom[  807] = 'h9ea315b4; 	    wvalid_rom[  807] = 0; 
    i_addr_rom[  808] = 'h00000794; 	    d_addr_rom[  808] = 'h00000d0c; 	    wdata_rom[  808] = 'h77af0c48; 	    wvalid_rom[  808] = 0; 
    i_addr_rom[  809] = 'h00000724; 	    d_addr_rom[  809] = 'h00000ce8; 	    wdata_rom[  809] = 'h3b9654fd; 	    wvalid_rom[  809] = 1; 
    i_addr_rom[  810] = 'h0000020c; 	    d_addr_rom[  810] = 'h00000970; 	    wdata_rom[  810] = 'h81265467; 	    wvalid_rom[  810] = 0; 
    i_addr_rom[  811] = 'h000005c0; 	    d_addr_rom[  811] = 'h00000820; 	    wdata_rom[  811] = 'h599da9b7; 	    wvalid_rom[  811] = 0; 
    i_addr_rom[  812] = 'h00000398; 	    d_addr_rom[  812] = 'h000008f4; 	    wdata_rom[  812] = 'h7b3e3627; 	    wvalid_rom[  812] = 0; 
    i_addr_rom[  813] = 'h0000010c; 	    d_addr_rom[  813] = 'h00000e64; 	    wdata_rom[  813] = 'h570e7d87; 	    wvalid_rom[  813] = 0; 
    i_addr_rom[  814] = 'h000004ac; 	    d_addr_rom[  814] = 'h00000de4; 	    wdata_rom[  814] = 'hf02828a0; 	    wvalid_rom[  814] = 1; 
    i_addr_rom[  815] = 'h00000298; 	    d_addr_rom[  815] = 'h00000b30; 	    wdata_rom[  815] = 'h2185c0a7; 	    wvalid_rom[  815] = 1; 
    i_addr_rom[  816] = 'h00000000; 	    d_addr_rom[  816] = 'h00000a10; 	    wdata_rom[  816] = 'hc7065675; 	    wvalid_rom[  816] = 0; 
    i_addr_rom[  817] = 'h00000010; 	    d_addr_rom[  817] = 'h00000ee4; 	    wdata_rom[  817] = 'h7d83c747; 	    wvalid_rom[  817] = 1; 
    i_addr_rom[  818] = 'h000001d0; 	    d_addr_rom[  818] = 'h0000089c; 	    wdata_rom[  818] = 'h8bbd4676; 	    wvalid_rom[  818] = 0; 
    i_addr_rom[  819] = 'h00000264; 	    d_addr_rom[  819] = 'h00000dec; 	    wdata_rom[  819] = 'hd477ad3b; 	    wvalid_rom[  819] = 1; 
    i_addr_rom[  820] = 'h0000042c; 	    d_addr_rom[  820] = 'h00000dfc; 	    wdata_rom[  820] = 'h3209e6c4; 	    wvalid_rom[  820] = 0; 
    i_addr_rom[  821] = 'h00000628; 	    d_addr_rom[  821] = 'h00000ee8; 	    wdata_rom[  821] = 'hdf51076b; 	    wvalid_rom[  821] = 1; 
    i_addr_rom[  822] = 'h000003c0; 	    d_addr_rom[  822] = 'h00000d94; 	    wdata_rom[  822] = 'hd66ed539; 	    wvalid_rom[  822] = 1; 
    i_addr_rom[  823] = 'h000003c4; 	    d_addr_rom[  823] = 'h00000d10; 	    wdata_rom[  823] = 'h5c60d4ca; 	    wvalid_rom[  823] = 0; 
    i_addr_rom[  824] = 'h00000170; 	    d_addr_rom[  824] = 'h00000ba8; 	    wdata_rom[  824] = 'h927cba5e; 	    wvalid_rom[  824] = 0; 
    i_addr_rom[  825] = 'h0000066c; 	    d_addr_rom[  825] = 'h00000d00; 	    wdata_rom[  825] = 'h2e859f3d; 	    wvalid_rom[  825] = 0; 
    i_addr_rom[  826] = 'h000001fc; 	    d_addr_rom[  826] = 'h00000d64; 	    wdata_rom[  826] = 'ha38a5af9; 	    wvalid_rom[  826] = 1; 
    i_addr_rom[  827] = 'h000001b8; 	    d_addr_rom[  827] = 'h00000df0; 	    wdata_rom[  827] = 'h41492e63; 	    wvalid_rom[  827] = 1; 
    i_addr_rom[  828] = 'h00000594; 	    d_addr_rom[  828] = 'h00000db8; 	    wdata_rom[  828] = 'hfd01934f; 	    wvalid_rom[  828] = 1; 
    i_addr_rom[  829] = 'h000003d0; 	    d_addr_rom[  829] = 'h00000ac8; 	    wdata_rom[  829] = 'h34c205e8; 	    wvalid_rom[  829] = 0; 
    i_addr_rom[  830] = 'h00000528; 	    d_addr_rom[  830] = 'h00000e60; 	    wdata_rom[  830] = 'hfe9d8a70; 	    wvalid_rom[  830] = 1; 
    i_addr_rom[  831] = 'h00000068; 	    d_addr_rom[  831] = 'h00000b3c; 	    wdata_rom[  831] = 'h20cdee65; 	    wvalid_rom[  831] = 1; 
    i_addr_rom[  832] = 'h000003b4; 	    d_addr_rom[  832] = 'h00000ccc; 	    wdata_rom[  832] = 'h7cb15dc3; 	    wvalid_rom[  832] = 1; 
    i_addr_rom[  833] = 'h00000250; 	    d_addr_rom[  833] = 'h00000a74; 	    wdata_rom[  833] = 'h06a4bbc6; 	    wvalid_rom[  833] = 0; 
    i_addr_rom[  834] = 'h000000dc; 	    d_addr_rom[  834] = 'h00000c00; 	    wdata_rom[  834] = 'he753c960; 	    wvalid_rom[  834] = 1; 
    i_addr_rom[  835] = 'h00000390; 	    d_addr_rom[  835] = 'h00000da0; 	    wdata_rom[  835] = 'h5855d8ce; 	    wvalid_rom[  835] = 1; 
    i_addr_rom[  836] = 'h000000bc; 	    d_addr_rom[  836] = 'h00000f10; 	    wdata_rom[  836] = 'hca972963; 	    wvalid_rom[  836] = 0; 
    i_addr_rom[  837] = 'h000000f0; 	    d_addr_rom[  837] = 'h000009ac; 	    wdata_rom[  837] = 'hdcceb029; 	    wvalid_rom[  837] = 1; 
    i_addr_rom[  838] = 'h0000048c; 	    d_addr_rom[  838] = 'h00000dec; 	    wdata_rom[  838] = 'h50a05050; 	    wvalid_rom[  838] = 0; 
    i_addr_rom[  839] = 'h000001a0; 	    d_addr_rom[  839] = 'h00000e00; 	    wdata_rom[  839] = 'h09202ac9; 	    wvalid_rom[  839] = 0; 
    i_addr_rom[  840] = 'h00000470; 	    d_addr_rom[  840] = 'h00000e7c; 	    wdata_rom[  840] = 'h10fc6395; 	    wvalid_rom[  840] = 1; 
    i_addr_rom[  841] = 'h00000174; 	    d_addr_rom[  841] = 'h00000e88; 	    wdata_rom[  841] = 'h4c13ae61; 	    wvalid_rom[  841] = 0; 
    i_addr_rom[  842] = 'h000007f8; 	    d_addr_rom[  842] = 'h0000089c; 	    wdata_rom[  842] = 'h587d1742; 	    wvalid_rom[  842] = 0; 
    i_addr_rom[  843] = 'h00000008; 	    d_addr_rom[  843] = 'h00000c3c; 	    wdata_rom[  843] = 'hddcffe9f; 	    wvalid_rom[  843] = 1; 
    i_addr_rom[  844] = 'h00000244; 	    d_addr_rom[  844] = 'h00000ee0; 	    wdata_rom[  844] = 'h534c5ac1; 	    wvalid_rom[  844] = 0; 
    i_addr_rom[  845] = 'h00000554; 	    d_addr_rom[  845] = 'h00000f98; 	    wdata_rom[  845] = 'hc457e5e6; 	    wvalid_rom[  845] = 1; 
    i_addr_rom[  846] = 'h00000624; 	    d_addr_rom[  846] = 'h00000e9c; 	    wdata_rom[  846] = 'h100946e3; 	    wvalid_rom[  846] = 1; 
    i_addr_rom[  847] = 'h000003e8; 	    d_addr_rom[  847] = 'h00000c18; 	    wdata_rom[  847] = 'ha8e2b0d9; 	    wvalid_rom[  847] = 1; 
    i_addr_rom[  848] = 'h00000670; 	    d_addr_rom[  848] = 'h00000e50; 	    wdata_rom[  848] = 'hd39ba74b; 	    wvalid_rom[  848] = 0; 
    i_addr_rom[  849] = 'h000007f8; 	    d_addr_rom[  849] = 'h00000c3c; 	    wdata_rom[  849] = 'hdb989979; 	    wvalid_rom[  849] = 0; 
    i_addr_rom[  850] = 'h00000134; 	    d_addr_rom[  850] = 'h00000a20; 	    wdata_rom[  850] = 'h41620df7; 	    wvalid_rom[  850] = 0; 
    i_addr_rom[  851] = 'h0000063c; 	    d_addr_rom[  851] = 'h00000b74; 	    wdata_rom[  851] = 'hf9712c2a; 	    wvalid_rom[  851] = 1; 
    i_addr_rom[  852] = 'h00000184; 	    d_addr_rom[  852] = 'h00000f64; 	    wdata_rom[  852] = 'h1e0dec51; 	    wvalid_rom[  852] = 0; 
    i_addr_rom[  853] = 'h000007a0; 	    d_addr_rom[  853] = 'h00000858; 	    wdata_rom[  853] = 'h320e1d27; 	    wvalid_rom[  853] = 1; 
    i_addr_rom[  854] = 'h000000b8; 	    d_addr_rom[  854] = 'h000009b0; 	    wdata_rom[  854] = 'hcf2e6961; 	    wvalid_rom[  854] = 0; 
    i_addr_rom[  855] = 'h00000298; 	    d_addr_rom[  855] = 'h00000ba4; 	    wdata_rom[  855] = 'h9aa15f20; 	    wvalid_rom[  855] = 1; 
    i_addr_rom[  856] = 'h00000314; 	    d_addr_rom[  856] = 'h000009b4; 	    wdata_rom[  856] = 'h18354c03; 	    wvalid_rom[  856] = 1; 
    i_addr_rom[  857] = 'h00000258; 	    d_addr_rom[  857] = 'h000009ac; 	    wdata_rom[  857] = 'h92f6c36c; 	    wvalid_rom[  857] = 0; 
    i_addr_rom[  858] = 'h000006fc; 	    d_addr_rom[  858] = 'h00000d78; 	    wdata_rom[  858] = 'ha18315ae; 	    wvalid_rom[  858] = 0; 
    i_addr_rom[  859] = 'h0000025c; 	    d_addr_rom[  859] = 'h00000a80; 	    wdata_rom[  859] = 'h20bd1dae; 	    wvalid_rom[  859] = 0; 
    i_addr_rom[  860] = 'h00000040; 	    d_addr_rom[  860] = 'h00000848; 	    wdata_rom[  860] = 'h22655e11; 	    wvalid_rom[  860] = 0; 
    i_addr_rom[  861] = 'h000001e4; 	    d_addr_rom[  861] = 'h00000ddc; 	    wdata_rom[  861] = 'h8a08fe98; 	    wvalid_rom[  861] = 0; 
    i_addr_rom[  862] = 'h000003f0; 	    d_addr_rom[  862] = 'h00000954; 	    wdata_rom[  862] = 'hb8f8e853; 	    wvalid_rom[  862] = 1; 
    i_addr_rom[  863] = 'h000006f4; 	    d_addr_rom[  863] = 'h00000a74; 	    wdata_rom[  863] = 'hf498f1cb; 	    wvalid_rom[  863] = 0; 
    i_addr_rom[  864] = 'h00000454; 	    d_addr_rom[  864] = 'h00000cb4; 	    wdata_rom[  864] = 'h57d43a8f; 	    wvalid_rom[  864] = 1; 
    i_addr_rom[  865] = 'h000005d8; 	    d_addr_rom[  865] = 'h00000fb4; 	    wdata_rom[  865] = 'h98244fb0; 	    wvalid_rom[  865] = 0; 
    i_addr_rom[  866] = 'h0000019c; 	    d_addr_rom[  866] = 'h00000a34; 	    wdata_rom[  866] = 'hffa906b1; 	    wvalid_rom[  866] = 0; 
    i_addr_rom[  867] = 'h000005f0; 	    d_addr_rom[  867] = 'h0000089c; 	    wdata_rom[  867] = 'hb4b58282; 	    wvalid_rom[  867] = 0; 
    i_addr_rom[  868] = 'h000001b4; 	    d_addr_rom[  868] = 'h00000dc8; 	    wdata_rom[  868] = 'h846a0348; 	    wvalid_rom[  868] = 1; 
    i_addr_rom[  869] = 'h00000590; 	    d_addr_rom[  869] = 'h00000e64; 	    wdata_rom[  869] = 'h169e9485; 	    wvalid_rom[  869] = 1; 
    i_addr_rom[  870] = 'h00000570; 	    d_addr_rom[  870] = 'h000008c4; 	    wdata_rom[  870] = 'h9fda57d8; 	    wvalid_rom[  870] = 0; 
    i_addr_rom[  871] = 'h00000350; 	    d_addr_rom[  871] = 'h00000df0; 	    wdata_rom[  871] = 'h6f50cd8e; 	    wvalid_rom[  871] = 1; 
    i_addr_rom[  872] = 'h000000dc; 	    d_addr_rom[  872] = 'h000008b0; 	    wdata_rom[  872] = 'h7f58a57b; 	    wvalid_rom[  872] = 1; 
    i_addr_rom[  873] = 'h00000568; 	    d_addr_rom[  873] = 'h00000918; 	    wdata_rom[  873] = 'h0a425225; 	    wvalid_rom[  873] = 1; 
    i_addr_rom[  874] = 'h00000774; 	    d_addr_rom[  874] = 'h00000ecc; 	    wdata_rom[  874] = 'heffe67db; 	    wvalid_rom[  874] = 0; 
    i_addr_rom[  875] = 'h0000041c; 	    d_addr_rom[  875] = 'h000009e4; 	    wdata_rom[  875] = 'h0414b8b1; 	    wvalid_rom[  875] = 1; 
    i_addr_rom[  876] = 'h0000031c; 	    d_addr_rom[  876] = 'h00000c70; 	    wdata_rom[  876] = 'h6adf73fd; 	    wvalid_rom[  876] = 0; 
    i_addr_rom[  877] = 'h00000554; 	    d_addr_rom[  877] = 'h00000ab4; 	    wdata_rom[  877] = 'ha6bdae29; 	    wvalid_rom[  877] = 1; 
    i_addr_rom[  878] = 'h000005c8; 	    d_addr_rom[  878] = 'h00000a14; 	    wdata_rom[  878] = 'h0f3c384d; 	    wvalid_rom[  878] = 0; 
    i_addr_rom[  879] = 'h00000140; 	    d_addr_rom[  879] = 'h00000f18; 	    wdata_rom[  879] = 'h3583e45b; 	    wvalid_rom[  879] = 1; 
    i_addr_rom[  880] = 'h00000160; 	    d_addr_rom[  880] = 'h00000d98; 	    wdata_rom[  880] = 'h8f3576e8; 	    wvalid_rom[  880] = 0; 
    i_addr_rom[  881] = 'h0000005c; 	    d_addr_rom[  881] = 'h00000f70; 	    wdata_rom[  881] = 'h08cc82e9; 	    wvalid_rom[  881] = 1; 
    i_addr_rom[  882] = 'h000005c4; 	    d_addr_rom[  882] = 'h00000dd8; 	    wdata_rom[  882] = 'h159eef9d; 	    wvalid_rom[  882] = 0; 
    i_addr_rom[  883] = 'h000001b0; 	    d_addr_rom[  883] = 'h00000b94; 	    wdata_rom[  883] = 'h172d4bdc; 	    wvalid_rom[  883] = 0; 
    i_addr_rom[  884] = 'h00000570; 	    d_addr_rom[  884] = 'h00000ef8; 	    wdata_rom[  884] = 'h27ab6dad; 	    wvalid_rom[  884] = 1; 
    i_addr_rom[  885] = 'h000003ac; 	    d_addr_rom[  885] = 'h00000f70; 	    wdata_rom[  885] = 'h902be43e; 	    wvalid_rom[  885] = 1; 
    i_addr_rom[  886] = 'h00000090; 	    d_addr_rom[  886] = 'h00000cb0; 	    wdata_rom[  886] = 'h546ee685; 	    wvalid_rom[  886] = 0; 
    i_addr_rom[  887] = 'h0000068c; 	    d_addr_rom[  887] = 'h00000dec; 	    wdata_rom[  887] = 'h4834ec4a; 	    wvalid_rom[  887] = 1; 
    i_addr_rom[  888] = 'h00000570; 	    d_addr_rom[  888] = 'h0000084c; 	    wdata_rom[  888] = 'hef980850; 	    wvalid_rom[  888] = 0; 
    i_addr_rom[  889] = 'h000000cc; 	    d_addr_rom[  889] = 'h00000d74; 	    wdata_rom[  889] = 'hebbec54e; 	    wvalid_rom[  889] = 1; 
    i_addr_rom[  890] = 'h0000007c; 	    d_addr_rom[  890] = 'h00000fcc; 	    wdata_rom[  890] = 'h86fee6ff; 	    wvalid_rom[  890] = 0; 
    i_addr_rom[  891] = 'h000000c0; 	    d_addr_rom[  891] = 'h00000be4; 	    wdata_rom[  891] = 'hcef45ed9; 	    wvalid_rom[  891] = 0; 
    i_addr_rom[  892] = 'h00000314; 	    d_addr_rom[  892] = 'h00000f60; 	    wdata_rom[  892] = 'he41d42d7; 	    wvalid_rom[  892] = 1; 
    i_addr_rom[  893] = 'h000000a8; 	    d_addr_rom[  893] = 'h00000d80; 	    wdata_rom[  893] = 'he34f3762; 	    wvalid_rom[  893] = 1; 
    i_addr_rom[  894] = 'h00000584; 	    d_addr_rom[  894] = 'h00000a60; 	    wdata_rom[  894] = 'h7707c3b7; 	    wvalid_rom[  894] = 0; 
    i_addr_rom[  895] = 'h000006f0; 	    d_addr_rom[  895] = 'h00000a10; 	    wdata_rom[  895] = 'h08a6aafa; 	    wvalid_rom[  895] = 1; 
    i_addr_rom[  896] = 'h00000700; 	    d_addr_rom[  896] = 'h00000c14; 	    wdata_rom[  896] = 'h033ad8c5; 	    wvalid_rom[  896] = 1; 
    i_addr_rom[  897] = 'h0000049c; 	    d_addr_rom[  897] = 'h00000ac4; 	    wdata_rom[  897] = 'h39e10b7a; 	    wvalid_rom[  897] = 1; 
    i_addr_rom[  898] = 'h000006c8; 	    d_addr_rom[  898] = 'h000008f0; 	    wdata_rom[  898] = 'h0c5fa1ce; 	    wvalid_rom[  898] = 0; 
    i_addr_rom[  899] = 'h00000184; 	    d_addr_rom[  899] = 'h00000cd8; 	    wdata_rom[  899] = 'h00cdf922; 	    wvalid_rom[  899] = 1; 
    i_addr_rom[  900] = 'h00000738; 	    d_addr_rom[  900] = 'h00000854; 	    wdata_rom[  900] = 'h2fa31440; 	    wvalid_rom[  900] = 0; 
    i_addr_rom[  901] = 'h00000240; 	    d_addr_rom[  901] = 'h00000c90; 	    wdata_rom[  901] = 'h4a4756b0; 	    wvalid_rom[  901] = 0; 
    i_addr_rom[  902] = 'h000006c0; 	    d_addr_rom[  902] = 'h00000910; 	    wdata_rom[  902] = 'h24533bfb; 	    wvalid_rom[  902] = 1; 
    i_addr_rom[  903] = 'h00000520; 	    d_addr_rom[  903] = 'h00000abc; 	    wdata_rom[  903] = 'hbcb19f80; 	    wvalid_rom[  903] = 1; 
    i_addr_rom[  904] = 'h00000080; 	    d_addr_rom[  904] = 'h00000e2c; 	    wdata_rom[  904] = 'hbb031292; 	    wvalid_rom[  904] = 0; 
    i_addr_rom[  905] = 'h0000014c; 	    d_addr_rom[  905] = 'h00000b34; 	    wdata_rom[  905] = 'hbcf3f7a2; 	    wvalid_rom[  905] = 1; 
    i_addr_rom[  906] = 'h00000230; 	    d_addr_rom[  906] = 'h00000a14; 	    wdata_rom[  906] = 'hf72309f2; 	    wvalid_rom[  906] = 0; 
    i_addr_rom[  907] = 'h0000070c; 	    d_addr_rom[  907] = 'h00000b64; 	    wdata_rom[  907] = 'hcb04ee59; 	    wvalid_rom[  907] = 0; 
    i_addr_rom[  908] = 'h0000046c; 	    d_addr_rom[  908] = 'h00000d4c; 	    wdata_rom[  908] = 'h8f70af37; 	    wvalid_rom[  908] = 1; 
    i_addr_rom[  909] = 'h000001b8; 	    d_addr_rom[  909] = 'h0000092c; 	    wdata_rom[  909] = 'hbb6e3a2c; 	    wvalid_rom[  909] = 0; 
    i_addr_rom[  910] = 'h000001dc; 	    d_addr_rom[  910] = 'h00000804; 	    wdata_rom[  910] = 'ha84069f6; 	    wvalid_rom[  910] = 0; 
    i_addr_rom[  911] = 'h000001e8; 	    d_addr_rom[  911] = 'h00000ddc; 	    wdata_rom[  911] = 'h9b891503; 	    wvalid_rom[  911] = 0; 
    i_addr_rom[  912] = 'h000007f8; 	    d_addr_rom[  912] = 'h00000d9c; 	    wdata_rom[  912] = 'h8ec3bb38; 	    wvalid_rom[  912] = 1; 
    i_addr_rom[  913] = 'h000002cc; 	    d_addr_rom[  913] = 'h00000db8; 	    wdata_rom[  913] = 'h55e37d8c; 	    wvalid_rom[  913] = 1; 
    i_addr_rom[  914] = 'h00000164; 	    d_addr_rom[  914] = 'h00000f18; 	    wdata_rom[  914] = 'hbdd7e22f; 	    wvalid_rom[  914] = 0; 
    i_addr_rom[  915] = 'h00000688; 	    d_addr_rom[  915] = 'h00000c58; 	    wdata_rom[  915] = 'h91ca8855; 	    wvalid_rom[  915] = 1; 
    i_addr_rom[  916] = 'h000006a4; 	    d_addr_rom[  916] = 'h00000950; 	    wdata_rom[  916] = 'h63b949c6; 	    wvalid_rom[  916] = 1; 
    i_addr_rom[  917] = 'h00000090; 	    d_addr_rom[  917] = 'h000009a8; 	    wdata_rom[  917] = 'h775dcabb; 	    wvalid_rom[  917] = 0; 
    i_addr_rom[  918] = 'h00000464; 	    d_addr_rom[  918] = 'h00000f9c; 	    wdata_rom[  918] = 'hd170d03d; 	    wvalid_rom[  918] = 1; 
    i_addr_rom[  919] = 'h00000740; 	    d_addr_rom[  919] = 'h00000a1c; 	    wdata_rom[  919] = 'hb8f486da; 	    wvalid_rom[  919] = 1; 
    i_addr_rom[  920] = 'h00000118; 	    d_addr_rom[  920] = 'h00000df0; 	    wdata_rom[  920] = 'h9d819a55; 	    wvalid_rom[  920] = 0; 
    i_addr_rom[  921] = 'h00000564; 	    d_addr_rom[  921] = 'h00000efc; 	    wdata_rom[  921] = 'h54e4312a; 	    wvalid_rom[  921] = 0; 
    i_addr_rom[  922] = 'h0000065c; 	    d_addr_rom[  922] = 'h00000d04; 	    wdata_rom[  922] = 'h4f6afc4b; 	    wvalid_rom[  922] = 1; 
    i_addr_rom[  923] = 'h000006d0; 	    d_addr_rom[  923] = 'h00000e04; 	    wdata_rom[  923] = 'hb3d5f3c0; 	    wvalid_rom[  923] = 0; 
    i_addr_rom[  924] = 'h00000798; 	    d_addr_rom[  924] = 'h00000c88; 	    wdata_rom[  924] = 'hba8b6d2b; 	    wvalid_rom[  924] = 0; 
    i_addr_rom[  925] = 'h00000378; 	    d_addr_rom[  925] = 'h00000c4c; 	    wdata_rom[  925] = 'h7a93d4a1; 	    wvalid_rom[  925] = 0; 
    i_addr_rom[  926] = 'h000005d0; 	    d_addr_rom[  926] = 'h00000f24; 	    wdata_rom[  926] = 'h0a312de9; 	    wvalid_rom[  926] = 1; 
    i_addr_rom[  927] = 'h00000358; 	    d_addr_rom[  927] = 'h00000d30; 	    wdata_rom[  927] = 'hf19a3d4a; 	    wvalid_rom[  927] = 0; 
    i_addr_rom[  928] = 'h00000678; 	    d_addr_rom[  928] = 'h00000f28; 	    wdata_rom[  928] = 'h45ccd706; 	    wvalid_rom[  928] = 1; 
    i_addr_rom[  929] = 'h000004a8; 	    d_addr_rom[  929] = 'h000009e8; 	    wdata_rom[  929] = 'hb259c942; 	    wvalid_rom[  929] = 0; 
    i_addr_rom[  930] = 'h000005bc; 	    d_addr_rom[  930] = 'h00000bdc; 	    wdata_rom[  930] = 'h4dc9f2b4; 	    wvalid_rom[  930] = 1; 
    i_addr_rom[  931] = 'h00000214; 	    d_addr_rom[  931] = 'h00000e9c; 	    wdata_rom[  931] = 'heb2b2f3b; 	    wvalid_rom[  931] = 1; 
    i_addr_rom[  932] = 'h000003f8; 	    d_addr_rom[  932] = 'h00000df0; 	    wdata_rom[  932] = 'he20f75d4; 	    wvalid_rom[  932] = 0; 
    i_addr_rom[  933] = 'h00000714; 	    d_addr_rom[  933] = 'h00000c2c; 	    wdata_rom[  933] = 'he49ad786; 	    wvalid_rom[  933] = 1; 
    i_addr_rom[  934] = 'h00000114; 	    d_addr_rom[  934] = 'h00000bb8; 	    wdata_rom[  934] = 'h47948766; 	    wvalid_rom[  934] = 1; 
    i_addr_rom[  935] = 'h00000190; 	    d_addr_rom[  935] = 'h00000eb4; 	    wdata_rom[  935] = 'he5de0076; 	    wvalid_rom[  935] = 1; 
    i_addr_rom[  936] = 'h0000027c; 	    d_addr_rom[  936] = 'h000008b0; 	    wdata_rom[  936] = 'h1f5e9a5e; 	    wvalid_rom[  936] = 1; 
    i_addr_rom[  937] = 'h000001c4; 	    d_addr_rom[  937] = 'h0000081c; 	    wdata_rom[  937] = 'h7ebc0249; 	    wvalid_rom[  937] = 1; 
    i_addr_rom[  938] = 'h00000230; 	    d_addr_rom[  938] = 'h00000f8c; 	    wdata_rom[  938] = 'h9037e787; 	    wvalid_rom[  938] = 0; 
    i_addr_rom[  939] = 'h000001d0; 	    d_addr_rom[  939] = 'h0000083c; 	    wdata_rom[  939] = 'hbe5fe24a; 	    wvalid_rom[  939] = 1; 
    i_addr_rom[  940] = 'h00000030; 	    d_addr_rom[  940] = 'h00000894; 	    wdata_rom[  940] = 'he2f17f0c; 	    wvalid_rom[  940] = 1; 
    i_addr_rom[  941] = 'h00000154; 	    d_addr_rom[  941] = 'h00000844; 	    wdata_rom[  941] = 'h92f96fe0; 	    wvalid_rom[  941] = 1; 
    i_addr_rom[  942] = 'h000005ec; 	    d_addr_rom[  942] = 'h00000f50; 	    wdata_rom[  942] = 'h2278949b; 	    wvalid_rom[  942] = 0; 
    i_addr_rom[  943] = 'h0000059c; 	    d_addr_rom[  943] = 'h000008ec; 	    wdata_rom[  943] = 'hc6159490; 	    wvalid_rom[  943] = 0; 
    i_addr_rom[  944] = 'h00000490; 	    d_addr_rom[  944] = 'h00000f44; 	    wdata_rom[  944] = 'h1d0e8c03; 	    wvalid_rom[  944] = 0; 
    i_addr_rom[  945] = 'h000005bc; 	    d_addr_rom[  945] = 'h00000b18; 	    wdata_rom[  945] = 'h95a9b41a; 	    wvalid_rom[  945] = 1; 
    i_addr_rom[  946] = 'h00000374; 	    d_addr_rom[  946] = 'h00000b58; 	    wdata_rom[  946] = 'h114fd842; 	    wvalid_rom[  946] = 1; 
    i_addr_rom[  947] = 'h000006ac; 	    d_addr_rom[  947] = 'h00000ff4; 	    wdata_rom[  947] = 'hd5d3f896; 	    wvalid_rom[  947] = 0; 
    i_addr_rom[  948] = 'h00000414; 	    d_addr_rom[  948] = 'h00000a2c; 	    wdata_rom[  948] = 'h371663df; 	    wvalid_rom[  948] = 1; 
    i_addr_rom[  949] = 'h000001d8; 	    d_addr_rom[  949] = 'h00000a28; 	    wdata_rom[  949] = 'h80f00181; 	    wvalid_rom[  949] = 1; 
    i_addr_rom[  950] = 'h00000080; 	    d_addr_rom[  950] = 'h00000b5c; 	    wdata_rom[  950] = 'hbd919d67; 	    wvalid_rom[  950] = 1; 
    i_addr_rom[  951] = 'h000007a8; 	    d_addr_rom[  951] = 'h00000e14; 	    wdata_rom[  951] = 'he36507a7; 	    wvalid_rom[  951] = 0; 
    i_addr_rom[  952] = 'h000007f8; 	    d_addr_rom[  952] = 'h00000f88; 	    wdata_rom[  952] = 'h41c41997; 	    wvalid_rom[  952] = 0; 
    i_addr_rom[  953] = 'h00000054; 	    d_addr_rom[  953] = 'h0000098c; 	    wdata_rom[  953] = 'h8ee2f91c; 	    wvalid_rom[  953] = 1; 
    i_addr_rom[  954] = 'h000004f0; 	    d_addr_rom[  954] = 'h00000998; 	    wdata_rom[  954] = 'h7820a2fb; 	    wvalid_rom[  954] = 0; 
    i_addr_rom[  955] = 'h000005a0; 	    d_addr_rom[  955] = 'h000009a8; 	    wdata_rom[  955] = 'h17d645b9; 	    wvalid_rom[  955] = 0; 
    i_addr_rom[  956] = 'h000002fc; 	    d_addr_rom[  956] = 'h00000dd4; 	    wdata_rom[  956] = 'h8d5cb6f9; 	    wvalid_rom[  956] = 0; 
    i_addr_rom[  957] = 'h00000188; 	    d_addr_rom[  957] = 'h00000b4c; 	    wdata_rom[  957] = 'h913c11d5; 	    wvalid_rom[  957] = 0; 
    i_addr_rom[  958] = 'h00000260; 	    d_addr_rom[  958] = 'h00000e24; 	    wdata_rom[  958] = 'hdf180506; 	    wvalid_rom[  958] = 0; 
    i_addr_rom[  959] = 'h000004a8; 	    d_addr_rom[  959] = 'h00000ab4; 	    wdata_rom[  959] = 'hd8be3527; 	    wvalid_rom[  959] = 1; 
    i_addr_rom[  960] = 'h00000250; 	    d_addr_rom[  960] = 'h00000b88; 	    wdata_rom[  960] = 'h58aeddb7; 	    wvalid_rom[  960] = 1; 
    i_addr_rom[  961] = 'h0000075c; 	    d_addr_rom[  961] = 'h00000928; 	    wdata_rom[  961] = 'h89f05b4f; 	    wvalid_rom[  961] = 0; 
    i_addr_rom[  962] = 'h00000640; 	    d_addr_rom[  962] = 'h00000e80; 	    wdata_rom[  962] = 'hf41f156c; 	    wvalid_rom[  962] = 0; 
    i_addr_rom[  963] = 'h000007f0; 	    d_addr_rom[  963] = 'h00000e30; 	    wdata_rom[  963] = 'hddd7dcb5; 	    wvalid_rom[  963] = 0; 
    i_addr_rom[  964] = 'h000002c4; 	    d_addr_rom[  964] = 'h00000e74; 	    wdata_rom[  964] = 'hd95e95f5; 	    wvalid_rom[  964] = 0; 
    i_addr_rom[  965] = 'h0000048c; 	    d_addr_rom[  965] = 'h00000c88; 	    wdata_rom[  965] = 'h6a89fe26; 	    wvalid_rom[  965] = 1; 
    i_addr_rom[  966] = 'h000004e8; 	    d_addr_rom[  966] = 'h00000ff0; 	    wdata_rom[  966] = 'h7f5b816f; 	    wvalid_rom[  966] = 0; 
    i_addr_rom[  967] = 'h000001dc; 	    d_addr_rom[  967] = 'h00000a88; 	    wdata_rom[  967] = 'h1f4b2ec0; 	    wvalid_rom[  967] = 1; 
    i_addr_rom[  968] = 'h000007f8; 	    d_addr_rom[  968] = 'h00000cf4; 	    wdata_rom[  968] = 'h1125f1af; 	    wvalid_rom[  968] = 1; 
    i_addr_rom[  969] = 'h000005c4; 	    d_addr_rom[  969] = 'h00000e34; 	    wdata_rom[  969] = 'h7ebf27fb; 	    wvalid_rom[  969] = 1; 
    i_addr_rom[  970] = 'h000000e0; 	    d_addr_rom[  970] = 'h00000970; 	    wdata_rom[  970] = 'h7778bda2; 	    wvalid_rom[  970] = 1; 
    i_addr_rom[  971] = 'h000007b0; 	    d_addr_rom[  971] = 'h00000e8c; 	    wdata_rom[  971] = 'h9159afc0; 	    wvalid_rom[  971] = 0; 
    i_addr_rom[  972] = 'h00000078; 	    d_addr_rom[  972] = 'h00000bb8; 	    wdata_rom[  972] = 'h0798d639; 	    wvalid_rom[  972] = 0; 
    i_addr_rom[  973] = 'h0000057c; 	    d_addr_rom[  973] = 'h00000d9c; 	    wdata_rom[  973] = 'hf2feb175; 	    wvalid_rom[  973] = 0; 
    i_addr_rom[  974] = 'h0000068c; 	    d_addr_rom[  974] = 'h00000dcc; 	    wdata_rom[  974] = 'h38de805c; 	    wvalid_rom[  974] = 0; 
    i_addr_rom[  975] = 'h00000390; 	    d_addr_rom[  975] = 'h00000f2c; 	    wdata_rom[  975] = 'h0d1b7f27; 	    wvalid_rom[  975] = 1; 
    i_addr_rom[  976] = 'h00000690; 	    d_addr_rom[  976] = 'h00000ffc; 	    wdata_rom[  976] = 'hd1c24e78; 	    wvalid_rom[  976] = 1; 
    i_addr_rom[  977] = 'h000000c0; 	    d_addr_rom[  977] = 'h00000820; 	    wdata_rom[  977] = 'he140a22b; 	    wvalid_rom[  977] = 0; 
    i_addr_rom[  978] = 'h00000340; 	    d_addr_rom[  978] = 'h00000e34; 	    wdata_rom[  978] = 'ha3b4bf55; 	    wvalid_rom[  978] = 1; 
    i_addr_rom[  979] = 'h0000054c; 	    d_addr_rom[  979] = 'h00000c88; 	    wdata_rom[  979] = 'hfc9bffb1; 	    wvalid_rom[  979] = 0; 
    i_addr_rom[  980] = 'h000007f0; 	    d_addr_rom[  980] = 'h00000e2c; 	    wdata_rom[  980] = 'h7a8be436; 	    wvalid_rom[  980] = 0; 
    i_addr_rom[  981] = 'h000002a0; 	    d_addr_rom[  981] = 'h00000d1c; 	    wdata_rom[  981] = 'hbf51474c; 	    wvalid_rom[  981] = 1; 
    i_addr_rom[  982] = 'h0000076c; 	    d_addr_rom[  982] = 'h000008cc; 	    wdata_rom[  982] = 'h3b4e9a62; 	    wvalid_rom[  982] = 0; 
    i_addr_rom[  983] = 'h00000320; 	    d_addr_rom[  983] = 'h00000d10; 	    wdata_rom[  983] = 'h10c784ca; 	    wvalid_rom[  983] = 0; 
    i_addr_rom[  984] = 'h000007a0; 	    d_addr_rom[  984] = 'h00000964; 	    wdata_rom[  984] = 'heb799e7f; 	    wvalid_rom[  984] = 1; 
    i_addr_rom[  985] = 'h0000008c; 	    d_addr_rom[  985] = 'h00000ff8; 	    wdata_rom[  985] = 'hf472ddc0; 	    wvalid_rom[  985] = 0; 
    i_addr_rom[  986] = 'h000000e0; 	    d_addr_rom[  986] = 'h00000edc; 	    wdata_rom[  986] = 'h756c3951; 	    wvalid_rom[  986] = 0; 
    i_addr_rom[  987] = 'h000006d8; 	    d_addr_rom[  987] = 'h00000b6c; 	    wdata_rom[  987] = 'hb662a083; 	    wvalid_rom[  987] = 0; 
    i_addr_rom[  988] = 'h00000304; 	    d_addr_rom[  988] = 'h00000844; 	    wdata_rom[  988] = 'h3c46b74a; 	    wvalid_rom[  988] = 1; 
    i_addr_rom[  989] = 'h00000364; 	    d_addr_rom[  989] = 'h00000d3c; 	    wdata_rom[  989] = 'hcf833908; 	    wvalid_rom[  989] = 0; 
    i_addr_rom[  990] = 'h000003dc; 	    d_addr_rom[  990] = 'h00000a18; 	    wdata_rom[  990] = 'h17f9bc9c; 	    wvalid_rom[  990] = 1; 
    i_addr_rom[  991] = 'h00000188; 	    d_addr_rom[  991] = 'h00000a90; 	    wdata_rom[  991] = 'h3047cf5d; 	    wvalid_rom[  991] = 1; 
    i_addr_rom[  992] = 'h00000258; 	    d_addr_rom[  992] = 'h00000dfc; 	    wdata_rom[  992] = 'h9a5c108a; 	    wvalid_rom[  992] = 0; 
    i_addr_rom[  993] = 'h00000324; 	    d_addr_rom[  993] = 'h00000d34; 	    wdata_rom[  993] = 'h0ac6f30b; 	    wvalid_rom[  993] = 1; 
    i_addr_rom[  994] = 'h000003e4; 	    d_addr_rom[  994] = 'h00000c44; 	    wdata_rom[  994] = 'hcb3db475; 	    wvalid_rom[  994] = 1; 
    i_addr_rom[  995] = 'h00000204; 	    d_addr_rom[  995] = 'h000009ac; 	    wdata_rom[  995] = 'h78816803; 	    wvalid_rom[  995] = 0; 
    i_addr_rom[  996] = 'h00000320; 	    d_addr_rom[  996] = 'h00000d3c; 	    wdata_rom[  996] = 'h671313b5; 	    wvalid_rom[  996] = 0; 
    i_addr_rom[  997] = 'h000000bc; 	    d_addr_rom[  997] = 'h00000e40; 	    wdata_rom[  997] = 'hd5fad3e5; 	    wvalid_rom[  997] = 1; 
    i_addr_rom[  998] = 'h0000002c; 	    d_addr_rom[  998] = 'h00000e7c; 	    wdata_rom[  998] = 'h0ab7ed28; 	    wvalid_rom[  998] = 1; 
    i_addr_rom[  999] = 'h00000608; 	    d_addr_rom[  999] = 'h00000f2c; 	    wdata_rom[  999] = 'he45319a2; 	    wvalid_rom[  999] = 0; 
    i_addr_rom[ 1000] = 'h000004d4; 	    d_addr_rom[ 1000] = 'h000009b8; 	    wdata_rom[ 1000] = 'h3cb2af9f; 	    wvalid_rom[ 1000] = 0; 
    i_addr_rom[ 1001] = 'h000004cc; 	    d_addr_rom[ 1001] = 'h00000c40; 	    wdata_rom[ 1001] = 'hc748b69c; 	    wvalid_rom[ 1001] = 1; 
    i_addr_rom[ 1002] = 'h00000798; 	    d_addr_rom[ 1002] = 'h00000bd4; 	    wdata_rom[ 1002] = 'h63b9e388; 	    wvalid_rom[ 1002] = 0; 
    i_addr_rom[ 1003] = 'h00000048; 	    d_addr_rom[ 1003] = 'h00000c84; 	    wdata_rom[ 1003] = 'ha7a24ab5; 	    wvalid_rom[ 1003] = 0; 
    i_addr_rom[ 1004] = 'h0000002c; 	    d_addr_rom[ 1004] = 'h00000ed4; 	    wdata_rom[ 1004] = 'h1e3bf8db; 	    wvalid_rom[ 1004] = 1; 
    i_addr_rom[ 1005] = 'h0000034c; 	    d_addr_rom[ 1005] = 'h00000f8c; 	    wdata_rom[ 1005] = 'h4b14670d; 	    wvalid_rom[ 1005] = 1; 
    i_addr_rom[ 1006] = 'h00000640; 	    d_addr_rom[ 1006] = 'h00000ba0; 	    wdata_rom[ 1006] = 'hda550a0e; 	    wvalid_rom[ 1006] = 1; 
    i_addr_rom[ 1007] = 'h0000036c; 	    d_addr_rom[ 1007] = 'h00000df8; 	    wdata_rom[ 1007] = 'h81a652d5; 	    wvalid_rom[ 1007] = 1; 
    i_addr_rom[ 1008] = 'h00000734; 	    d_addr_rom[ 1008] = 'h00000c3c; 	    wdata_rom[ 1008] = 'h501b3732; 	    wvalid_rom[ 1008] = 1; 
    i_addr_rom[ 1009] = 'h000003c0; 	    d_addr_rom[ 1009] = 'h00000d68; 	    wdata_rom[ 1009] = 'h2d94a4ff; 	    wvalid_rom[ 1009] = 1; 
    i_addr_rom[ 1010] = 'h000004a4; 	    d_addr_rom[ 1010] = 'h00000f1c; 	    wdata_rom[ 1010] = 'h70b2ee72; 	    wvalid_rom[ 1010] = 1; 
    i_addr_rom[ 1011] = 'h00000624; 	    d_addr_rom[ 1011] = 'h00000dac; 	    wdata_rom[ 1011] = 'hff2e3a37; 	    wvalid_rom[ 1011] = 1; 
    i_addr_rom[ 1012] = 'h00000094; 	    d_addr_rom[ 1012] = 'h00000948; 	    wdata_rom[ 1012] = 'haab062e9; 	    wvalid_rom[ 1012] = 1; 
    i_addr_rom[ 1013] = 'h00000190; 	    d_addr_rom[ 1013] = 'h00000c6c; 	    wdata_rom[ 1013] = 'h8d18643c; 	    wvalid_rom[ 1013] = 1; 
    i_addr_rom[ 1014] = 'h000002f4; 	    d_addr_rom[ 1014] = 'h00000be8; 	    wdata_rom[ 1014] = 'h067abc72; 	    wvalid_rom[ 1014] = 1; 
    i_addr_rom[ 1015] = 'h000003f0; 	    d_addr_rom[ 1015] = 'h00000c64; 	    wdata_rom[ 1015] = 'h90aaba51; 	    wvalid_rom[ 1015] = 0; 
    i_addr_rom[ 1016] = 'h0000053c; 	    d_addr_rom[ 1016] = 'h00000af0; 	    wdata_rom[ 1016] = 'h216194a2; 	    wvalid_rom[ 1016] = 0; 
    i_addr_rom[ 1017] = 'h00000504; 	    d_addr_rom[ 1017] = 'h000008fc; 	    wdata_rom[ 1017] = 'h79573836; 	    wvalid_rom[ 1017] = 0; 
    i_addr_rom[ 1018] = 'h00000620; 	    d_addr_rom[ 1018] = 'h00000ab4; 	    wdata_rom[ 1018] = 'h2d781b13; 	    wvalid_rom[ 1018] = 1; 
    i_addr_rom[ 1019] = 'h00000430; 	    d_addr_rom[ 1019] = 'h00000f0c; 	    wdata_rom[ 1019] = 'h27f8b8df; 	    wvalid_rom[ 1019] = 0; 
    i_addr_rom[ 1020] = 'h00000558; 	    d_addr_rom[ 1020] = 'h00000c38; 	    wdata_rom[ 1020] = 'hd53e299d; 	    wvalid_rom[ 1020] = 0; 
    i_addr_rom[ 1021] = 'h00000234; 	    d_addr_rom[ 1021] = 'h00000b74; 	    wdata_rom[ 1021] = 'h5951ca12; 	    wvalid_rom[ 1021] = 1; 
    i_addr_rom[ 1022] = 'h0000068c; 	    d_addr_rom[ 1022] = 'h00000e94; 	    wdata_rom[ 1022] = 'h61110d96; 	    wvalid_rom[ 1022] = 1; 
    i_addr_rom[ 1023] = 'h0000078c; 	    d_addr_rom[ 1023] = 'h00000844; 	    wdata_rom[ 1023] = 'ha5fb4cd1; 	    wvalid_rom[ 1023] = 0; 

end
// for icache 
wire            i_rvalid_pipe;
wire            i_rready_pipe;
wire    [31:0]  i_raddr_pipe;
wire    [31:0]  i_rdata_pipe;
wire            i_rvalid;
wire            i_rready;
// icache && arbiter 
wire    [31:0]  i_raddr;
wire    [31:0]  i_rdata;
wire            i_rlast;
wire    [2:0]   i_rsize;
wire    [7:0]   i_rlen;
// icache_debug
reg             i_rvalid_ff;
reg     [31:0]  i_raddr_ff;
reg             i_error_reg;
reg             i_pass_reg;
wire    [31:0]  i_correct_data;

// for dcache
wire    [31:0]  d_addr_pipe;
wire            d_rvalid_pipe;
wire            d_rready_pipe;
wire    [31:0]  d_rdata_pipe;
wire            d_wvalid_pipe;
wire            d_wready_pipe;
wire    [31:0]  d_wdata_pipe;
wire    [3:0]   d_wstrb_pipe;
// dcache && arbiter
wire            d_rvalid;
wire            d_rready;
wire    [31:0]  d_raddr;
wire    [31:0]  d_rdata;
wire            d_rlast;
wire    [2:0]   d_rsize;
wire    [7:0]   d_rlen;
wire            d_wvalid;
wire            d_wready;
wire    [31:0]  d_waddr;
wire    [31:0]  d_wdata;
wire    [3:0]   d_wstrb;
wire            d_wlast;
wire    [2:0]   d_wsize;
wire    [7:0]   d_wlen;
wire            d_bvalid;
wire            d_bready;
// dcache_debug
reg             d_rvalid_ff;
reg             d_wvalid_ff;
reg     [31:0]  d_wdata_ff;
reg     [31:0]  d_addr_ff;
reg             d_error_reg;
reg             d_pass_reg;
wire    [31:0]  d_correct_data;

// arbiter with main mem
wire    [31:0]  araddr;
wire            arvalid;
wire            arready;
wire    [7:0]   arlen;
wire    [2:0]   arsize;
wire    [1:0]   arburst;
wire    [31:0]  rdata;
wire    [1:0]   rresp;
wire            rvalid;
wire            rready;
wire            rlast;
wire    [31:0]  awaddr;
wire            awvalid;
wire            awready;
wire    [7:0]   awlen;
wire    [2:0]   awsize;
wire    [1:0]   awburst;
wire    [31:0]  wdata;
wire    [3:0]   wstrb;
wire            wvalid;
wire            wready;
wire            wlast;
wire    [1:0]   bresp;
wire            bvalid;
wire            bready;

assign i_raddr_pipe = i_addr_rom[i_test_index];
assign i_correct_data = data_ram[i_raddr_ff >> 2];
assign i_rvalid_pipe = 1'b1;
// simulate IF1-IF2 register i_rvalid_ff && i_raddr_ff
always @(posedge clk) begin
    if(!rstn) begin
        i_rvalid_ff <= 0;
        i_raddr_ff <= 0;
    end
    else if(!(i_rvalid_ff && !i_rready_pipe))begin
        i_rvalid_ff <= i_rvalid_pipe;
        i_raddr_ff <= i_raddr_pipe;
    end
end
// update i_test_index
always @(posedge clk) begin
    if(!rstn) begin
        i_test_index <= 0;
        i_pass_reg <= 0;
    end
    else if (i_test_index >= (TOTAL_WORD_NUM / 2-1)) begin
        i_test_index <= (TOTAL_WORD_NUM / 2-1);
        i_pass_reg <= 1;
    end
    else if(!(i_rvalid_ff && !i_rready_pipe) && !i_error_reg) begin
        i_test_index <= i_test_index + 1;
    end
end
// update i_error 
always @(posedge clk) begin
    if(!rstn) begin
        i_error_reg <= 0;
    end
    else if(i_error_reg) begin
        i_error_reg <= 1;
    end
    else if(i_rvalid_ff && i_rready_pipe) begin
        i_error_reg <= !(i_rdata_pipe  == i_correct_data);
    end
end

assign d_addr_pipe           = d_addr_rom[d_test_index];
assign d_correct_data   = data_ram[d_addr_ff >> 2];
assign d_rvalid_pipe         = !wvalid_rom[d_test_index];
assign d_wvalid_pipe         = wvalid_rom[d_test_index];
assign d_wdata_pipe          = wdata_rom[d_test_index];
assign d_wstrb_pipe          = d_wvalid_pipe ? 4'b1111 : 4'b0000;
// simulate EX-MEM register
always @(posedge clk) begin
    if(!rstn) begin
        d_rvalid_ff <= 0;
        d_addr_ff   <= 0;
        d_wvalid_ff <= 0;
        d_wdata_ff  <= 0;
    end
    else if(!(d_rvalid_ff && !d_rready_pipe) && !(d_wvalid_ff && !d_wready_pipe))begin
        d_rvalid_ff <= d_rvalid_pipe;
        d_addr_ff   <= d_addr_pipe;
        d_wvalid_ff <= d_wvalid_pipe;
        d_wdata_ff  <= d_wdata_pipe;
    end
end
// update d_test_index
always @(posedge clk) begin
    if(!rstn) begin
        d_test_index    <= TOTAL_WORD_NUM / 2;
        d_pass_reg      <= 0;
    end
    else if (d_test_index >= (TOTAL_WORD_NUM-1)) begin
        d_test_index    <= (TOTAL_WORD_NUM-1);
        d_pass_reg      <= 1;
    end
    else if(!(d_rvalid_ff && !d_rready_pipe)  && !(d_wvalid_ff && !d_wready_pipe) && !d_error_reg) begin
        d_test_index    <= d_test_index + 1;
    end
end
// update data_ram
always @(posedge clk) begin
    if(d_wvalid_ff && d_wready_pipe) begin
        data_ram[d_addr_ff >> 2] <= d_wdata_ff;
    end
end
// update d_error 
always @(posedge clk) begin
    if(!rstn) begin
        d_error_reg <= 0;
    end
    else if(d_error_reg) begin
        d_error_reg <= 1;
    end
    else if(d_rvalid_ff && d_rready_pipe) begin
        d_error_reg <= !(d_rdata_pipe  == d_correct_data);
    end
end

    wire mem_icache_dataOK, mem_dcache_dataOK;
    wire icache_mem_req, dcache_mem_req;
    wire [127:0] dout_mem_icache, dout_mem_dcache;

Icache #(
  .index_width          (INDEX_WIDTH),
  .offset_width    (WORD_OFFSET_WIDTH)
)
icache_dut (
    .clk      (clk ),
    .rstn     (rstn ),
    .test1    (),
    .test2    (),
    .test3    (),
    // .rvalid   (i_rvalid_pipe ),
    // .rready   (i_rready_pipe ),
    // .raddr    (i_raddr_pipe ),
    // .rdata    (i_rdata_pipe ),

    // .i_rvalid (i_rvalid ),
    // .i_rready (i_rready ),
    // .i_raddr  (i_raddr ),
    // .i_rdata  (i_rdata ),
    // .i_rlast  (i_rlast ),
    // .i_rsize  (i_rsize ),
    // .i_rlen   (i_rlen)
    .addr_pipeline_icache    (i_raddr_pipe),
    .dout_icache_pipeline   (i_rdata_pipe),
    .flag_icache_pipeline   (),
    .pipeline_icache_valid  (i_rvalid_pipe),
    .icache_pipeline_ready  (i_rready_pipe),

    .pipeline_icache_opcode (0),
    .pipeline_icache_opflag (1'b0),
    .pipeline_icache_ctrl   (0),
    .icache_pipeline_stall  (),
    
    //l1-axi
    .addr_icache_mem        (i_raddr),
    .din_mem_icache         (dout_mem_icache),
    
    .icache_mem_req         (icache_mem_req),
    .icache_mem_size        (i_rsize),

    // .mem_icache_addrOK      (),
    .mem_icache_dataOK      (mem_icache_dataOK)
);

ReturnBuffer#(
    .offset_width(WORD_OFFSET_WIDTH)
)
icache_returnbuf(
    .clk                (clk),
    .rstn               (rstn),
    .cache_mem_req      (icache_mem_req),
    .mem_cache_dataOK   (mem_icache_dataOK),
    .dout_mem_cache     (dout_mem_icache),
    .rready             (i_rready),
    .rdata              (i_rdata),
    .rlast              (i_rlast)
);

    wire    wr_type;
    wire    [2:0]dcache_mem_size;
    wire    dcache_pipeline_ready;
    wire    type_pipeline_dcache;
    wire    [31:0]addr_dcache_mem;

    assign d_raddr=addr_dcache_mem;
    assign d_waddr=addr_dcache_mem;

    assign d_rsize=dcache_mem_size;
    assign d_wsize=dcache_mem_size;
    assign d_rvalid=wr_type?0:dcache_mem_req;
    assign d_wvalid=wr_type?dcache_mem_req:0;

    assign d_rready=dcache_pipeline_ready;
    assign d_wready=dcache_pipeline_ready;

    assign type_pipeline_dcache=d_rvalid_pipe?0:d_wvalid_pipe;

Dcache #(
    .index_width        (INDEX_WIDTH ),
    .offset_width  (WORD_OFFSET_WIDTH )
)
dcache_dut (
    // .clk      (clk ),
    // .rstn     (rstn ),
    // .addr     (d_addr_pipe ),
    // .rvalid   (d_rvalid_pipe ),
    // .rready   (d_rready_pipe ),
    // .rdata    (d_rdata_pipe ),
    // .wvalid   (d_wvalid_pipe ),
    // .wready   (d_wready_pipe ),
    // .wdata    (d_wdata_pipe ),
    // .wstrb    (d_wstrb_pipe ),
    // .d_rvalid (d_rvalid ),
    // .d_rready (d_rready ),
    // .d_raddr  (d_raddr ),
    // .d_rdata  (d_rdata ),
    // .d_rlast  (d_rlast ),
    // .d_rsize  (d_rsize ),
    // .d_rlen   (d_rlen ),
    // .d_wvalid (d_wvalid ),
    // .d_wready (d_wready ),
    // .d_waddr  (d_waddr ),
    // .d_wdata  (d_wdata ),
    // .d_wstrb  (d_wstrb ),
    // .d_wlast  (d_wlast ),
    // .d_wsize  (d_wsize ),
    // .d_wlen   (d_wlen ),
    // .d_bvalid (d_bvalid ),
    // .d_bready (d_bready )
    
    .clk                    (clk),
    .rstn                   (rstn),
    .test1                  (),
    .test2                  (),
    .test3                  (),

    .addr_pipeline_dcache   (d_addr_pipe),
    .din_pipeline_dcache    (d_wdata_pipe),
    .dout_dcache_pipeline   (d_rdata_pipe),
    .type_pipeline_dcache   (type_pipeline_dcache),

    .pipeline_dcache_valid  (d_rvalid_pipe&d_wvalid_pipe),
    .dcache_pipeline_ready  (dcache_pipeline_ready),

    .pipeline_dcache_wstrb  (d_wstrb_pipe),
    .pipeline_dcache_opcode (0),
    .pipeline_dcache_opflag (1'b0),
    .pipeline_dcache_ctrl   (0),
    .dcache_pipeline_stall  (),

    .addr_dcache_mem        (addr_dcache_mem),
    .dout_dcache_mem        (d_wdata),
    .din_mem_dcache         (dout_mem_dcache),

    .dcache_mem_req         (dcache_mem_req),
    .dcache_mem_wr          (wr_type),
    .dcache_mem_size        (dcache_mem_size),
    .dcache_mem_wstrb       (d_wstrb),
    // .mem_dcache_addrOK      (),
    .mem_dcache_dataOK      (mem_dcache_dataOK)
);

ReturnBuffer#(
    .offset_width(WORD_OFFSET_WIDTH)
)
dcache_returnbuf(
    .clk                (clk),
    .rstn               (rstn),
    .cache_mem_req      (dcache_mem_req),
    .mem_cache_dataOK   (mem_dcache_dataOK),
    .dout_mem_cache     (dout_mem_dcache),
    .rready             (d_rready),
    .rdata              (d_rdata),
    .rlast              (d_rlast)
);


axi_arbiter axi_arbiter_dut (
    .clk      (clk ),
    .rstn     (rstn ),
    .i_rvalid (i_rvalid ),
    .i_rready (i_rready ),
    .i_raddr  (i_raddr ),
    .i_rdata  (i_rdata ),
    .i_rlast  (i_rlast ),
    .i_rsize  (i_rsize ),
    .i_rlen   (1 ),
    .d_rvalid (d_rvalid ),
    .d_rready (d_rready ),
    .d_raddr  (d_raddr ),
    .d_rdata  (d_rdata ),
    .d_rlast  (d_rlast ),
    .d_rsize  (d_rsize ),
    .d_rlen   (d_rlen ),
    .d_wvalid (d_wvalid ),
    .d_wready (d_wready ),
    .d_waddr  (d_waddr ),
    .d_wdata  (d_wdata ),
    .d_wstrb  (d_wstrb ),
    .d_wlast  (d_wlast ),
    .d_wsize  (d_wsize ),
    .d_wlen   (d_wlen ),
    .d_bvalid (d_bvalid ),
    .d_bready (d_bready ),
    .araddr   (araddr ),
    .arvalid  (arvalid ),
    .arready  (arready ),
    .arlen    (arlen ),
    .arsize   (arsize ),
    .arburst  (arburst ),
    .rdata    (rdata ),
    .rresp    (rresp ),
    .rvalid   (rvalid ),
    .rready   (rready ),
    .rlast    (rlast ),
    .awaddr   (awaddr ),
    .awvalid  (awvalid ),
    .awready  (awready ),
    .awlen    (awlen ),
    .awsize   (awsize ),
    .awburst  (awburst ),
    .wdata    (wdata ),
    .wstrb    (wstrb ),
    .wvalid   (wvalid ),
    .wready   (wready ),
    .wlast    (wlast ),
    .bresp    (bresp ),
    .bvalid   (bvalid ),
    .bready   (bready)
);
main_memory main_mem(
    .s_aclk         (clk ),
    .s_aresetn      (rstn ),
    .s_axi_araddr   (araddr ),
    .s_axi_arburst  (arburst ),
    .s_axi_arid     (4'b0),
    .s_axi_arlen    (arlen ),
    .s_axi_arready  (arready ),
    .s_axi_arsize   (arsize ),
    .s_axi_arvalid  (arvalid ),
    .s_axi_awaddr   (awaddr ),
    .s_axi_awburst  (awburst ),
    .s_axi_awid     (4'b0),
    .s_axi_awlen    (awlen ),
    .s_axi_awready  (awready ),
    .s_axi_awsize   (awsize ),
    .s_axi_awvalid  (awvalid ),
    .s_axi_bid      (),
    .s_axi_bready   (bready ),
    .s_axi_bresp    (bresp ),
    .s_axi_bvalid   (bvalid ),
    .s_axi_rdata    (rdata ),
    .s_axi_rid      (),
    .s_axi_rlast    (rlast ),
    .s_axi_rready   (rready ),
    .s_axi_rresp    (rresp ),
    .s_axi_rvalid   (rvalid ),
    .s_axi_wdata    (wdata ),
    .s_axi_wlast    (wlast ),
    .s_axi_wready   (wready ),
    .s_axi_wstrb    (wstrb ),
    .s_axi_wvalid   (wvalid )
);
endmodule
