module IPCP_pre(



);

localparam  = ;

endmodule