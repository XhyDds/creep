module fetch_buffer_v2 (
    input [31:0]pc,
    input clk,rstn,flush,stall,
    input if0,if1,icache_valid,
    input [1:0]plv,
    input [63:0]irin,
    input [63:0]pre,
    // input [63:0]
    input flag,
    input [15:0]excp_arg,
    //flag==1表示2个有效，flag==0表示1个有效
    //[0:31]为pc小，0-后一条指令（[63:32]）无效 1-有效
    output [31:0]ir0,ir1,pc0,pc1,
    output stall_fetch_buffer,valid0,valid1,
    output [1:0]plv0,plv1,
    output [63:0]pre0,pre1,
    output [15:0]excp_arg0,excp_arg1
);
    reg [31:0]buffer[0:15];//15为0，14最新，0最旧，是否会溢出？
    reg [31:0]bufferpc[0:15];
    reg [66:0]pre_and_valid_and_plv[0:15];
    reg [15:0]excp_arg[0:15];
    reg [3:0]pointer;//0~15
    wire [31:0]ir[0:1];
    assign ir[0]=irin[31:0];
    assign ir[1]=irin[63:32];
    assign ir0=buffer[pointer==15?pointer:pointer+1];
    assign ir1=buffer[pointer];
    assign pc0=bufferpc[pointer==15?pointer:pointer+1];
    assign pc1=bufferpc[pointer];
    assign stall_fetch_buffer=(pointer<=1);
    assign valid0=pre_and_valid_and_plv[pointer==15?pointer:pointer+1][2];
    assign valid1=pre_and_valid_and_plv[pointer][2];
    assign plv0=pre_and_valid_and_plv[pointer==15?pointer:pointer+1][1:0];
    assign plv1=pre_and_valid_and_plv[pointer][1:0];
    assign pre0=pre_and_valid_and_plv[pointer==15?pointer:pointer+1][66:3];
    assign pre1=pre_and_valid_and_plv[pointer][66:3];
    assign excp_arg0=excp_arg[pointer==15?pointer:pointer+1];
    assign excp_arg1=excp_arg[pointer];
    wire [3:0]flag4p=icache_valid?(flag?4'b0010:4'b0001):4'b0000;
    wire [3:0]flag4=icache_valid?(flag?4'b0001:4'b0000):4'b1111;
    wire [3:0]flag4m=icache_valid?(flag?4'b0000:4'b1111):4'b1110;

    always @(posedge clk,negedge rstn) begin
        if(!rstn|flush) 
            begin
                pointer<=15;
                for (i=0;i<16;i=i+1) begin
                        buffer[i]<=0;
                        bufferpc[i]<=0;
                        pre_and_valid_and_plv[i]<=0;
                end
            end
        else if(!stall)
            begin
                if(icache_valid)
                    if (flag) 
                        begin
                            genvar i;
                            generate for(i = 0 ; i < 13; i = i + 1) begin : U
                                buffer[i]<=buffer[i+2];
                                bufferpc[i]<=bufferpc[i+2];
                                pre_and_valid_and_plv[i]<=pre_and_valid_and_plv[i+2];
                                excp_arg[i]<=excp_arg[i+2];
                            end
                            endgenerate
                            buffer[13]<=ir[0];
                            bufferpc[13]<=pc;
                            pre_and_valid_and_plv[13]<={pre,1'b1,plv};
                            excp_arg[13]<=excp_arg;
                            buffer[14]<=ir[1];
                            bufferpc[14]<=pc+4;
                            pre_and_valid_and_plv[14]<={pre,1'b1,plv};
                            excp_arg[14]<=0;
                        end
                    else 
                        begin
                            genvar i;
                            generate for(i = 0 ; i < 14; i = i + 1) begin : U
                                buffer[i]<=buffer[i+1];
                                bufferpc[i]<=bufferpc[i+1];
                                pre_and_valid_and_plv[i]<=pre_and_valid_and_plv[i+1];
                                excp_arg[i]<=excp_arg[i+1];
                            end
                            endgenerate
                            buffer[14]<=ir[0];
                            bufferpc[14]<=pc;
                            pre_and_valid_and_plv[14]<={pre,1'b1,plv};
                            excp_arg[14]<=excp_arg;
                        end
                if(if1)
                    if(if0) pointer<=(pointer==14|pointer==15)?(15-flag4p):(pointer-flag4m);//取两个
                    else pointer<=(pointer==15)?(15-flag4p):(pointer-flag4);//取一个
                else
                    pointer<=pointer-flag4p;
                //有下面走，上面不走的情况吗？
            end
    end
endmodule
