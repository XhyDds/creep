//hash函数for单输入
module single_hash#(
    parameter DATA_width=32,
    parameter HASH_width=32
) (
    input [DATA_width-1:0] data_raw,
    output[HASH_width-1:0] data_hashed
);
    
endmodule