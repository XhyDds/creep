module inst_pre#(

)(

);
endmodule